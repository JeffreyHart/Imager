magic
tech scmos
timestamp 1354157810
<< ntransistor >>
rect 18 879 21 881
rect 32 872 34 875
rect 63 879 66 881
rect 77 872 79 875
rect 13 862 15 865
rect 23 862 25 865
rect 108 879 111 881
rect 122 872 124 875
rect 58 862 60 865
rect 68 862 70 865
rect 153 879 156 881
rect 167 872 169 875
rect 103 862 105 865
rect 113 862 115 865
rect 198 879 201 881
rect 212 872 214 875
rect 148 862 150 865
rect 158 862 160 865
rect 243 879 246 881
rect 257 872 259 875
rect 193 862 195 865
rect 203 862 205 865
rect 288 879 291 881
rect 302 872 304 875
rect 238 862 240 865
rect 248 862 250 865
rect 333 879 336 881
rect 347 872 349 875
rect 283 862 285 865
rect 293 862 295 865
rect 378 879 381 881
rect 392 872 394 875
rect 328 862 330 865
rect 338 862 340 865
rect 423 879 426 881
rect 437 872 439 875
rect 373 862 375 865
rect 383 862 385 865
rect 468 879 471 881
rect 482 872 484 875
rect 418 862 420 865
rect 428 862 430 865
rect 513 879 516 881
rect 527 872 529 875
rect 463 862 465 865
rect 473 862 475 865
rect 558 879 561 881
rect 572 872 574 875
rect 508 862 510 865
rect 518 862 520 865
rect 603 879 606 881
rect 617 872 619 875
rect 553 862 555 865
rect 563 862 565 865
rect 648 879 651 881
rect 662 872 664 875
rect 598 862 600 865
rect 608 862 610 865
rect 693 879 696 881
rect 707 872 709 875
rect 643 862 645 865
rect 653 862 655 865
rect 738 879 741 881
rect 752 872 754 875
rect 688 862 690 865
rect 698 862 700 865
rect 783 879 786 881
rect 797 872 799 875
rect 733 862 735 865
rect 743 862 745 865
rect 828 879 831 881
rect 842 872 844 875
rect 778 862 780 865
rect 788 862 790 865
rect 873 879 876 881
rect 887 872 889 875
rect 823 862 825 865
rect 833 862 835 865
rect 868 862 870 865
rect 878 862 880 865
rect 18 834 21 836
rect 32 827 34 830
rect 63 834 66 836
rect 77 827 79 830
rect 13 817 15 820
rect 23 817 25 820
rect 108 834 111 836
rect 122 827 124 830
rect 58 817 60 820
rect 68 817 70 820
rect 153 834 156 836
rect 167 827 169 830
rect 103 817 105 820
rect 113 817 115 820
rect 198 834 201 836
rect 212 827 214 830
rect 148 817 150 820
rect 158 817 160 820
rect 243 834 246 836
rect 257 827 259 830
rect 193 817 195 820
rect 203 817 205 820
rect 288 834 291 836
rect 302 827 304 830
rect 238 817 240 820
rect 248 817 250 820
rect 333 834 336 836
rect 347 827 349 830
rect 283 817 285 820
rect 293 817 295 820
rect 378 834 381 836
rect 392 827 394 830
rect 328 817 330 820
rect 338 817 340 820
rect 423 834 426 836
rect 437 827 439 830
rect 373 817 375 820
rect 383 817 385 820
rect 468 834 471 836
rect 482 827 484 830
rect 418 817 420 820
rect 428 817 430 820
rect 513 834 516 836
rect 527 827 529 830
rect 463 817 465 820
rect 473 817 475 820
rect 558 834 561 836
rect 572 827 574 830
rect 508 817 510 820
rect 518 817 520 820
rect 603 834 606 836
rect 617 827 619 830
rect 553 817 555 820
rect 563 817 565 820
rect 648 834 651 836
rect 662 827 664 830
rect 598 817 600 820
rect 608 817 610 820
rect 693 834 696 836
rect 707 827 709 830
rect 643 817 645 820
rect 653 817 655 820
rect 738 834 741 836
rect 752 827 754 830
rect 688 817 690 820
rect 698 817 700 820
rect 783 834 786 836
rect 797 827 799 830
rect 733 817 735 820
rect 743 817 745 820
rect 828 834 831 836
rect 842 827 844 830
rect 778 817 780 820
rect 788 817 790 820
rect 873 834 876 836
rect 887 827 889 830
rect 823 817 825 820
rect 833 817 835 820
rect 868 817 870 820
rect 878 817 880 820
rect 18 789 21 791
rect 32 782 34 785
rect 63 789 66 791
rect 77 782 79 785
rect 13 772 15 775
rect 23 772 25 775
rect 108 789 111 791
rect 122 782 124 785
rect 58 772 60 775
rect 68 772 70 775
rect 153 789 156 791
rect 167 782 169 785
rect 103 772 105 775
rect 113 772 115 775
rect 198 789 201 791
rect 212 782 214 785
rect 148 772 150 775
rect 158 772 160 775
rect 243 789 246 791
rect 257 782 259 785
rect 193 772 195 775
rect 203 772 205 775
rect 288 789 291 791
rect 302 782 304 785
rect 238 772 240 775
rect 248 772 250 775
rect 333 789 336 791
rect 347 782 349 785
rect 283 772 285 775
rect 293 772 295 775
rect 378 789 381 791
rect 392 782 394 785
rect 328 772 330 775
rect 338 772 340 775
rect 423 789 426 791
rect 437 782 439 785
rect 373 772 375 775
rect 383 772 385 775
rect 468 789 471 791
rect 482 782 484 785
rect 418 772 420 775
rect 428 772 430 775
rect 513 789 516 791
rect 527 782 529 785
rect 463 772 465 775
rect 473 772 475 775
rect 558 789 561 791
rect 572 782 574 785
rect 508 772 510 775
rect 518 772 520 775
rect 603 789 606 791
rect 617 782 619 785
rect 553 772 555 775
rect 563 772 565 775
rect 648 789 651 791
rect 662 782 664 785
rect 598 772 600 775
rect 608 772 610 775
rect 693 789 696 791
rect 707 782 709 785
rect 643 772 645 775
rect 653 772 655 775
rect 738 789 741 791
rect 752 782 754 785
rect 688 772 690 775
rect 698 772 700 775
rect 783 789 786 791
rect 797 782 799 785
rect 733 772 735 775
rect 743 772 745 775
rect 828 789 831 791
rect 842 782 844 785
rect 778 772 780 775
rect 788 772 790 775
rect 873 789 876 791
rect 887 782 889 785
rect 823 772 825 775
rect 833 772 835 775
rect 868 772 870 775
rect 878 772 880 775
rect 18 744 21 746
rect 32 737 34 740
rect 63 744 66 746
rect 77 737 79 740
rect 13 727 15 730
rect 23 727 25 730
rect 108 744 111 746
rect 122 737 124 740
rect 58 727 60 730
rect 68 727 70 730
rect 153 744 156 746
rect 167 737 169 740
rect 103 727 105 730
rect 113 727 115 730
rect 198 744 201 746
rect 212 737 214 740
rect 148 727 150 730
rect 158 727 160 730
rect 243 744 246 746
rect 257 737 259 740
rect 193 727 195 730
rect 203 727 205 730
rect 288 744 291 746
rect 302 737 304 740
rect 238 727 240 730
rect 248 727 250 730
rect 333 744 336 746
rect 347 737 349 740
rect 283 727 285 730
rect 293 727 295 730
rect 378 744 381 746
rect 392 737 394 740
rect 328 727 330 730
rect 338 727 340 730
rect 423 744 426 746
rect 437 737 439 740
rect 373 727 375 730
rect 383 727 385 730
rect 468 744 471 746
rect 482 737 484 740
rect 418 727 420 730
rect 428 727 430 730
rect 513 744 516 746
rect 527 737 529 740
rect 463 727 465 730
rect 473 727 475 730
rect 558 744 561 746
rect 572 737 574 740
rect 508 727 510 730
rect 518 727 520 730
rect 603 744 606 746
rect 617 737 619 740
rect 553 727 555 730
rect 563 727 565 730
rect 648 744 651 746
rect 662 737 664 740
rect 598 727 600 730
rect 608 727 610 730
rect 693 744 696 746
rect 707 737 709 740
rect 643 727 645 730
rect 653 727 655 730
rect 738 744 741 746
rect 752 737 754 740
rect 688 727 690 730
rect 698 727 700 730
rect 783 744 786 746
rect 797 737 799 740
rect 733 727 735 730
rect 743 727 745 730
rect 828 744 831 746
rect 842 737 844 740
rect 778 727 780 730
rect 788 727 790 730
rect 873 744 876 746
rect 887 737 889 740
rect 823 727 825 730
rect 833 727 835 730
rect 868 727 870 730
rect 878 727 880 730
rect 18 699 21 701
rect 32 692 34 695
rect 63 699 66 701
rect 77 692 79 695
rect 13 682 15 685
rect 23 682 25 685
rect 108 699 111 701
rect 122 692 124 695
rect 58 682 60 685
rect 68 682 70 685
rect 153 699 156 701
rect 167 692 169 695
rect 103 682 105 685
rect 113 682 115 685
rect 198 699 201 701
rect 212 692 214 695
rect 148 682 150 685
rect 158 682 160 685
rect 243 699 246 701
rect 257 692 259 695
rect 193 682 195 685
rect 203 682 205 685
rect 288 699 291 701
rect 302 692 304 695
rect 238 682 240 685
rect 248 682 250 685
rect 333 699 336 701
rect 347 692 349 695
rect 283 682 285 685
rect 293 682 295 685
rect 378 699 381 701
rect 392 692 394 695
rect 328 682 330 685
rect 338 682 340 685
rect 423 699 426 701
rect 437 692 439 695
rect 373 682 375 685
rect 383 682 385 685
rect 468 699 471 701
rect 482 692 484 695
rect 418 682 420 685
rect 428 682 430 685
rect 513 699 516 701
rect 527 692 529 695
rect 463 682 465 685
rect 473 682 475 685
rect 558 699 561 701
rect 572 692 574 695
rect 508 682 510 685
rect 518 682 520 685
rect 603 699 606 701
rect 617 692 619 695
rect 553 682 555 685
rect 563 682 565 685
rect 648 699 651 701
rect 662 692 664 695
rect 598 682 600 685
rect 608 682 610 685
rect 693 699 696 701
rect 707 692 709 695
rect 643 682 645 685
rect 653 682 655 685
rect 738 699 741 701
rect 752 692 754 695
rect 688 682 690 685
rect 698 682 700 685
rect 783 699 786 701
rect 797 692 799 695
rect 733 682 735 685
rect 743 682 745 685
rect 828 699 831 701
rect 842 692 844 695
rect 778 682 780 685
rect 788 682 790 685
rect 873 699 876 701
rect 887 692 889 695
rect 823 682 825 685
rect 833 682 835 685
rect 868 682 870 685
rect 878 682 880 685
rect 18 654 21 656
rect 32 647 34 650
rect 63 654 66 656
rect 77 647 79 650
rect 13 637 15 640
rect 23 637 25 640
rect 108 654 111 656
rect 122 647 124 650
rect 58 637 60 640
rect 68 637 70 640
rect 153 654 156 656
rect 167 647 169 650
rect 103 637 105 640
rect 113 637 115 640
rect 198 654 201 656
rect 212 647 214 650
rect 148 637 150 640
rect 158 637 160 640
rect 243 654 246 656
rect 257 647 259 650
rect 193 637 195 640
rect 203 637 205 640
rect 288 654 291 656
rect 302 647 304 650
rect 238 637 240 640
rect 248 637 250 640
rect 333 654 336 656
rect 347 647 349 650
rect 283 637 285 640
rect 293 637 295 640
rect 378 654 381 656
rect 392 647 394 650
rect 328 637 330 640
rect 338 637 340 640
rect 423 654 426 656
rect 437 647 439 650
rect 373 637 375 640
rect 383 637 385 640
rect 468 654 471 656
rect 482 647 484 650
rect 418 637 420 640
rect 428 637 430 640
rect 513 654 516 656
rect 527 647 529 650
rect 463 637 465 640
rect 473 637 475 640
rect 558 654 561 656
rect 572 647 574 650
rect 508 637 510 640
rect 518 637 520 640
rect 603 654 606 656
rect 617 647 619 650
rect 553 637 555 640
rect 563 637 565 640
rect 648 654 651 656
rect 662 647 664 650
rect 598 637 600 640
rect 608 637 610 640
rect 693 654 696 656
rect 707 647 709 650
rect 643 637 645 640
rect 653 637 655 640
rect 738 654 741 656
rect 752 647 754 650
rect 688 637 690 640
rect 698 637 700 640
rect 783 654 786 656
rect 797 647 799 650
rect 733 637 735 640
rect 743 637 745 640
rect 828 654 831 656
rect 842 647 844 650
rect 778 637 780 640
rect 788 637 790 640
rect 873 654 876 656
rect 887 647 889 650
rect 823 637 825 640
rect 833 637 835 640
rect 868 637 870 640
rect 878 637 880 640
rect 18 609 21 611
rect 32 602 34 605
rect 63 609 66 611
rect 77 602 79 605
rect 13 592 15 595
rect 23 592 25 595
rect 108 609 111 611
rect 122 602 124 605
rect 58 592 60 595
rect 68 592 70 595
rect 153 609 156 611
rect 167 602 169 605
rect 103 592 105 595
rect 113 592 115 595
rect 198 609 201 611
rect 212 602 214 605
rect 148 592 150 595
rect 158 592 160 595
rect 243 609 246 611
rect 257 602 259 605
rect 193 592 195 595
rect 203 592 205 595
rect 288 609 291 611
rect 302 602 304 605
rect 238 592 240 595
rect 248 592 250 595
rect 333 609 336 611
rect 347 602 349 605
rect 283 592 285 595
rect 293 592 295 595
rect 378 609 381 611
rect 392 602 394 605
rect 328 592 330 595
rect 338 592 340 595
rect 423 609 426 611
rect 437 602 439 605
rect 373 592 375 595
rect 383 592 385 595
rect 468 609 471 611
rect 482 602 484 605
rect 418 592 420 595
rect 428 592 430 595
rect 513 609 516 611
rect 527 602 529 605
rect 463 592 465 595
rect 473 592 475 595
rect 558 609 561 611
rect 572 602 574 605
rect 508 592 510 595
rect 518 592 520 595
rect 603 609 606 611
rect 617 602 619 605
rect 553 592 555 595
rect 563 592 565 595
rect 648 609 651 611
rect 662 602 664 605
rect 598 592 600 595
rect 608 592 610 595
rect 693 609 696 611
rect 707 602 709 605
rect 643 592 645 595
rect 653 592 655 595
rect 738 609 741 611
rect 752 602 754 605
rect 688 592 690 595
rect 698 592 700 595
rect 783 609 786 611
rect 797 602 799 605
rect 733 592 735 595
rect 743 592 745 595
rect 828 609 831 611
rect 842 602 844 605
rect 778 592 780 595
rect 788 592 790 595
rect 873 609 876 611
rect 887 602 889 605
rect 823 592 825 595
rect 833 592 835 595
rect 868 592 870 595
rect 878 592 880 595
rect 18 564 21 566
rect 32 557 34 560
rect 63 564 66 566
rect 77 557 79 560
rect 13 547 15 550
rect 23 547 25 550
rect 108 564 111 566
rect 122 557 124 560
rect 58 547 60 550
rect 68 547 70 550
rect 153 564 156 566
rect 167 557 169 560
rect 103 547 105 550
rect 113 547 115 550
rect 198 564 201 566
rect 212 557 214 560
rect 148 547 150 550
rect 158 547 160 550
rect 243 564 246 566
rect 257 557 259 560
rect 193 547 195 550
rect 203 547 205 550
rect 288 564 291 566
rect 302 557 304 560
rect 238 547 240 550
rect 248 547 250 550
rect 333 564 336 566
rect 347 557 349 560
rect 283 547 285 550
rect 293 547 295 550
rect 378 564 381 566
rect 392 557 394 560
rect 328 547 330 550
rect 338 547 340 550
rect 423 564 426 566
rect 437 557 439 560
rect 373 547 375 550
rect 383 547 385 550
rect 468 564 471 566
rect 482 557 484 560
rect 418 547 420 550
rect 428 547 430 550
rect 513 564 516 566
rect 527 557 529 560
rect 463 547 465 550
rect 473 547 475 550
rect 558 564 561 566
rect 572 557 574 560
rect 508 547 510 550
rect 518 547 520 550
rect 603 564 606 566
rect 617 557 619 560
rect 553 547 555 550
rect 563 547 565 550
rect 648 564 651 566
rect 662 557 664 560
rect 598 547 600 550
rect 608 547 610 550
rect 693 564 696 566
rect 707 557 709 560
rect 643 547 645 550
rect 653 547 655 550
rect 738 564 741 566
rect 752 557 754 560
rect 688 547 690 550
rect 698 547 700 550
rect 783 564 786 566
rect 797 557 799 560
rect 733 547 735 550
rect 743 547 745 550
rect 828 564 831 566
rect 842 557 844 560
rect 778 547 780 550
rect 788 547 790 550
rect 873 564 876 566
rect 887 557 889 560
rect 823 547 825 550
rect 833 547 835 550
rect 868 547 870 550
rect 878 547 880 550
rect 18 519 21 521
rect 32 512 34 515
rect 63 519 66 521
rect 77 512 79 515
rect 13 502 15 505
rect 23 502 25 505
rect 108 519 111 521
rect 122 512 124 515
rect 58 502 60 505
rect 68 502 70 505
rect 153 519 156 521
rect 167 512 169 515
rect 103 502 105 505
rect 113 502 115 505
rect 198 519 201 521
rect 212 512 214 515
rect 148 502 150 505
rect 158 502 160 505
rect 243 519 246 521
rect 257 512 259 515
rect 193 502 195 505
rect 203 502 205 505
rect 288 519 291 521
rect 302 512 304 515
rect 238 502 240 505
rect 248 502 250 505
rect 333 519 336 521
rect 347 512 349 515
rect 283 502 285 505
rect 293 502 295 505
rect 378 519 381 521
rect 392 512 394 515
rect 328 502 330 505
rect 338 502 340 505
rect 423 519 426 521
rect 437 512 439 515
rect 373 502 375 505
rect 383 502 385 505
rect 468 519 471 521
rect 482 512 484 515
rect 418 502 420 505
rect 428 502 430 505
rect 513 519 516 521
rect 527 512 529 515
rect 463 502 465 505
rect 473 502 475 505
rect 558 519 561 521
rect 572 512 574 515
rect 508 502 510 505
rect 518 502 520 505
rect 603 519 606 521
rect 617 512 619 515
rect 553 502 555 505
rect 563 502 565 505
rect 648 519 651 521
rect 662 512 664 515
rect 598 502 600 505
rect 608 502 610 505
rect 693 519 696 521
rect 707 512 709 515
rect 643 502 645 505
rect 653 502 655 505
rect 738 519 741 521
rect 752 512 754 515
rect 688 502 690 505
rect 698 502 700 505
rect 783 519 786 521
rect 797 512 799 515
rect 733 502 735 505
rect 743 502 745 505
rect 828 519 831 521
rect 842 512 844 515
rect 778 502 780 505
rect 788 502 790 505
rect 873 519 876 521
rect 887 512 889 515
rect 823 502 825 505
rect 833 502 835 505
rect 868 502 870 505
rect 878 502 880 505
rect 18 474 21 476
rect 32 467 34 470
rect 63 474 66 476
rect 77 467 79 470
rect 13 457 15 460
rect 23 457 25 460
rect 108 474 111 476
rect 122 467 124 470
rect 58 457 60 460
rect 68 457 70 460
rect 153 474 156 476
rect 167 467 169 470
rect 103 457 105 460
rect 113 457 115 460
rect 198 474 201 476
rect 212 467 214 470
rect 148 457 150 460
rect 158 457 160 460
rect 243 474 246 476
rect 257 467 259 470
rect 193 457 195 460
rect 203 457 205 460
rect 288 474 291 476
rect 302 467 304 470
rect 238 457 240 460
rect 248 457 250 460
rect 333 474 336 476
rect 347 467 349 470
rect 283 457 285 460
rect 293 457 295 460
rect 378 474 381 476
rect 392 467 394 470
rect 328 457 330 460
rect 338 457 340 460
rect 423 474 426 476
rect 437 467 439 470
rect 373 457 375 460
rect 383 457 385 460
rect 468 474 471 476
rect 482 467 484 470
rect 418 457 420 460
rect 428 457 430 460
rect 513 474 516 476
rect 527 467 529 470
rect 463 457 465 460
rect 473 457 475 460
rect 558 474 561 476
rect 572 467 574 470
rect 508 457 510 460
rect 518 457 520 460
rect 603 474 606 476
rect 617 467 619 470
rect 553 457 555 460
rect 563 457 565 460
rect 648 474 651 476
rect 662 467 664 470
rect 598 457 600 460
rect 608 457 610 460
rect 693 474 696 476
rect 707 467 709 470
rect 643 457 645 460
rect 653 457 655 460
rect 738 474 741 476
rect 752 467 754 470
rect 688 457 690 460
rect 698 457 700 460
rect 783 474 786 476
rect 797 467 799 470
rect 733 457 735 460
rect 743 457 745 460
rect 828 474 831 476
rect 842 467 844 470
rect 778 457 780 460
rect 788 457 790 460
rect 873 474 876 476
rect 887 467 889 470
rect 823 457 825 460
rect 833 457 835 460
rect 868 457 870 460
rect 878 457 880 460
rect 18 429 21 431
rect 32 422 34 425
rect 63 429 66 431
rect 77 422 79 425
rect 13 412 15 415
rect 23 412 25 415
rect 108 429 111 431
rect 122 422 124 425
rect 58 412 60 415
rect 68 412 70 415
rect 153 429 156 431
rect 167 422 169 425
rect 103 412 105 415
rect 113 412 115 415
rect 198 429 201 431
rect 212 422 214 425
rect 148 412 150 415
rect 158 412 160 415
rect 243 429 246 431
rect 257 422 259 425
rect 193 412 195 415
rect 203 412 205 415
rect 288 429 291 431
rect 302 422 304 425
rect 238 412 240 415
rect 248 412 250 415
rect 333 429 336 431
rect 347 422 349 425
rect 283 412 285 415
rect 293 412 295 415
rect 378 429 381 431
rect 392 422 394 425
rect 328 412 330 415
rect 338 412 340 415
rect 423 429 426 431
rect 437 422 439 425
rect 373 412 375 415
rect 383 412 385 415
rect 468 429 471 431
rect 482 422 484 425
rect 418 412 420 415
rect 428 412 430 415
rect 513 429 516 431
rect 527 422 529 425
rect 463 412 465 415
rect 473 412 475 415
rect 558 429 561 431
rect 572 422 574 425
rect 508 412 510 415
rect 518 412 520 415
rect 603 429 606 431
rect 617 422 619 425
rect 553 412 555 415
rect 563 412 565 415
rect 648 429 651 431
rect 662 422 664 425
rect 598 412 600 415
rect 608 412 610 415
rect 693 429 696 431
rect 707 422 709 425
rect 643 412 645 415
rect 653 412 655 415
rect 738 429 741 431
rect 752 422 754 425
rect 688 412 690 415
rect 698 412 700 415
rect 783 429 786 431
rect 797 422 799 425
rect 733 412 735 415
rect 743 412 745 415
rect 828 429 831 431
rect 842 422 844 425
rect 778 412 780 415
rect 788 412 790 415
rect 873 429 876 431
rect 887 422 889 425
rect 823 412 825 415
rect 833 412 835 415
rect 868 412 870 415
rect 878 412 880 415
rect 18 384 21 386
rect 32 377 34 380
rect 63 384 66 386
rect 77 377 79 380
rect 13 367 15 370
rect 23 367 25 370
rect 108 384 111 386
rect 122 377 124 380
rect 58 367 60 370
rect 68 367 70 370
rect 153 384 156 386
rect 167 377 169 380
rect 103 367 105 370
rect 113 367 115 370
rect 198 384 201 386
rect 212 377 214 380
rect 148 367 150 370
rect 158 367 160 370
rect 243 384 246 386
rect 257 377 259 380
rect 193 367 195 370
rect 203 367 205 370
rect 288 384 291 386
rect 302 377 304 380
rect 238 367 240 370
rect 248 367 250 370
rect 333 384 336 386
rect 347 377 349 380
rect 283 367 285 370
rect 293 367 295 370
rect 378 384 381 386
rect 392 377 394 380
rect 328 367 330 370
rect 338 367 340 370
rect 423 384 426 386
rect 437 377 439 380
rect 373 367 375 370
rect 383 367 385 370
rect 468 384 471 386
rect 482 377 484 380
rect 418 367 420 370
rect 428 367 430 370
rect 513 384 516 386
rect 527 377 529 380
rect 463 367 465 370
rect 473 367 475 370
rect 558 384 561 386
rect 572 377 574 380
rect 508 367 510 370
rect 518 367 520 370
rect 603 384 606 386
rect 617 377 619 380
rect 553 367 555 370
rect 563 367 565 370
rect 648 384 651 386
rect 662 377 664 380
rect 598 367 600 370
rect 608 367 610 370
rect 693 384 696 386
rect 707 377 709 380
rect 643 367 645 370
rect 653 367 655 370
rect 738 384 741 386
rect 752 377 754 380
rect 688 367 690 370
rect 698 367 700 370
rect 783 384 786 386
rect 797 377 799 380
rect 733 367 735 370
rect 743 367 745 370
rect 828 384 831 386
rect 842 377 844 380
rect 778 367 780 370
rect 788 367 790 370
rect 873 384 876 386
rect 887 377 889 380
rect 823 367 825 370
rect 833 367 835 370
rect 868 367 870 370
rect 878 367 880 370
rect 18 339 21 341
rect 32 332 34 335
rect 63 339 66 341
rect 77 332 79 335
rect 13 322 15 325
rect 23 322 25 325
rect 108 339 111 341
rect 122 332 124 335
rect 58 322 60 325
rect 68 322 70 325
rect 153 339 156 341
rect 167 332 169 335
rect 103 322 105 325
rect 113 322 115 325
rect 198 339 201 341
rect 212 332 214 335
rect 148 322 150 325
rect 158 322 160 325
rect 243 339 246 341
rect 257 332 259 335
rect 193 322 195 325
rect 203 322 205 325
rect 288 339 291 341
rect 302 332 304 335
rect 238 322 240 325
rect 248 322 250 325
rect 333 339 336 341
rect 347 332 349 335
rect 283 322 285 325
rect 293 322 295 325
rect 378 339 381 341
rect 392 332 394 335
rect 328 322 330 325
rect 338 322 340 325
rect 423 339 426 341
rect 437 332 439 335
rect 373 322 375 325
rect 383 322 385 325
rect 468 339 471 341
rect 482 332 484 335
rect 418 322 420 325
rect 428 322 430 325
rect 513 339 516 341
rect 527 332 529 335
rect 463 322 465 325
rect 473 322 475 325
rect 558 339 561 341
rect 572 332 574 335
rect 508 322 510 325
rect 518 322 520 325
rect 603 339 606 341
rect 617 332 619 335
rect 553 322 555 325
rect 563 322 565 325
rect 648 339 651 341
rect 662 332 664 335
rect 598 322 600 325
rect 608 322 610 325
rect 693 339 696 341
rect 707 332 709 335
rect 643 322 645 325
rect 653 322 655 325
rect 738 339 741 341
rect 752 332 754 335
rect 688 322 690 325
rect 698 322 700 325
rect 783 339 786 341
rect 797 332 799 335
rect 733 322 735 325
rect 743 322 745 325
rect 828 339 831 341
rect 842 332 844 335
rect 778 322 780 325
rect 788 322 790 325
rect 873 339 876 341
rect 887 332 889 335
rect 823 322 825 325
rect 833 322 835 325
rect 868 322 870 325
rect 878 322 880 325
rect 18 294 21 296
rect 32 287 34 290
rect 63 294 66 296
rect 77 287 79 290
rect 13 277 15 280
rect 23 277 25 280
rect 108 294 111 296
rect 122 287 124 290
rect 58 277 60 280
rect 68 277 70 280
rect 153 294 156 296
rect 167 287 169 290
rect 103 277 105 280
rect 113 277 115 280
rect 198 294 201 296
rect 212 287 214 290
rect 148 277 150 280
rect 158 277 160 280
rect 243 294 246 296
rect 257 287 259 290
rect 193 277 195 280
rect 203 277 205 280
rect 288 294 291 296
rect 302 287 304 290
rect 238 277 240 280
rect 248 277 250 280
rect 333 294 336 296
rect 347 287 349 290
rect 283 277 285 280
rect 293 277 295 280
rect 378 294 381 296
rect 392 287 394 290
rect 328 277 330 280
rect 338 277 340 280
rect 423 294 426 296
rect 437 287 439 290
rect 373 277 375 280
rect 383 277 385 280
rect 468 294 471 296
rect 482 287 484 290
rect 418 277 420 280
rect 428 277 430 280
rect 513 294 516 296
rect 527 287 529 290
rect 463 277 465 280
rect 473 277 475 280
rect 558 294 561 296
rect 572 287 574 290
rect 508 277 510 280
rect 518 277 520 280
rect 603 294 606 296
rect 617 287 619 290
rect 553 277 555 280
rect 563 277 565 280
rect 648 294 651 296
rect 662 287 664 290
rect 598 277 600 280
rect 608 277 610 280
rect 693 294 696 296
rect 707 287 709 290
rect 643 277 645 280
rect 653 277 655 280
rect 738 294 741 296
rect 752 287 754 290
rect 688 277 690 280
rect 698 277 700 280
rect 783 294 786 296
rect 797 287 799 290
rect 733 277 735 280
rect 743 277 745 280
rect 828 294 831 296
rect 842 287 844 290
rect 778 277 780 280
rect 788 277 790 280
rect 873 294 876 296
rect 887 287 889 290
rect 823 277 825 280
rect 833 277 835 280
rect 868 277 870 280
rect 878 277 880 280
rect 18 249 21 251
rect 32 242 34 245
rect 63 249 66 251
rect 77 242 79 245
rect 13 232 15 235
rect 23 232 25 235
rect 108 249 111 251
rect 122 242 124 245
rect 58 232 60 235
rect 68 232 70 235
rect 153 249 156 251
rect 167 242 169 245
rect 103 232 105 235
rect 113 232 115 235
rect 198 249 201 251
rect 212 242 214 245
rect 148 232 150 235
rect 158 232 160 235
rect 243 249 246 251
rect 257 242 259 245
rect 193 232 195 235
rect 203 232 205 235
rect 288 249 291 251
rect 302 242 304 245
rect 238 232 240 235
rect 248 232 250 235
rect 333 249 336 251
rect 347 242 349 245
rect 283 232 285 235
rect 293 232 295 235
rect 378 249 381 251
rect 392 242 394 245
rect 328 232 330 235
rect 338 232 340 235
rect 423 249 426 251
rect 437 242 439 245
rect 373 232 375 235
rect 383 232 385 235
rect 468 249 471 251
rect 482 242 484 245
rect 418 232 420 235
rect 428 232 430 235
rect 513 249 516 251
rect 527 242 529 245
rect 463 232 465 235
rect 473 232 475 235
rect 558 249 561 251
rect 572 242 574 245
rect 508 232 510 235
rect 518 232 520 235
rect 603 249 606 251
rect 617 242 619 245
rect 553 232 555 235
rect 563 232 565 235
rect 648 249 651 251
rect 662 242 664 245
rect 598 232 600 235
rect 608 232 610 235
rect 693 249 696 251
rect 707 242 709 245
rect 643 232 645 235
rect 653 232 655 235
rect 738 249 741 251
rect 752 242 754 245
rect 688 232 690 235
rect 698 232 700 235
rect 783 249 786 251
rect 797 242 799 245
rect 733 232 735 235
rect 743 232 745 235
rect 828 249 831 251
rect 842 242 844 245
rect 778 232 780 235
rect 788 232 790 235
rect 873 249 876 251
rect 887 242 889 245
rect 823 232 825 235
rect 833 232 835 235
rect 868 232 870 235
rect 878 232 880 235
rect 18 204 21 206
rect 32 197 34 200
rect 63 204 66 206
rect 77 197 79 200
rect 13 187 15 190
rect 23 187 25 190
rect 108 204 111 206
rect 122 197 124 200
rect 58 187 60 190
rect 68 187 70 190
rect 153 204 156 206
rect 167 197 169 200
rect 103 187 105 190
rect 113 187 115 190
rect 198 204 201 206
rect 212 197 214 200
rect 148 187 150 190
rect 158 187 160 190
rect 243 204 246 206
rect 257 197 259 200
rect 193 187 195 190
rect 203 187 205 190
rect 288 204 291 206
rect 302 197 304 200
rect 238 187 240 190
rect 248 187 250 190
rect 333 204 336 206
rect 347 197 349 200
rect 283 187 285 190
rect 293 187 295 190
rect 378 204 381 206
rect 392 197 394 200
rect 328 187 330 190
rect 338 187 340 190
rect 423 204 426 206
rect 437 197 439 200
rect 373 187 375 190
rect 383 187 385 190
rect 468 204 471 206
rect 482 197 484 200
rect 418 187 420 190
rect 428 187 430 190
rect 513 204 516 206
rect 527 197 529 200
rect 463 187 465 190
rect 473 187 475 190
rect 558 204 561 206
rect 572 197 574 200
rect 508 187 510 190
rect 518 187 520 190
rect 603 204 606 206
rect 617 197 619 200
rect 553 187 555 190
rect 563 187 565 190
rect 648 204 651 206
rect 662 197 664 200
rect 598 187 600 190
rect 608 187 610 190
rect 693 204 696 206
rect 707 197 709 200
rect 643 187 645 190
rect 653 187 655 190
rect 738 204 741 206
rect 752 197 754 200
rect 688 187 690 190
rect 698 187 700 190
rect 783 204 786 206
rect 797 197 799 200
rect 733 187 735 190
rect 743 187 745 190
rect 828 204 831 206
rect 842 197 844 200
rect 778 187 780 190
rect 788 187 790 190
rect 873 204 876 206
rect 887 197 889 200
rect 823 187 825 190
rect 833 187 835 190
rect 868 187 870 190
rect 878 187 880 190
rect 18 159 21 161
rect 32 152 34 155
rect 63 159 66 161
rect 77 152 79 155
rect 13 142 15 145
rect 23 142 25 145
rect 108 159 111 161
rect 122 152 124 155
rect 58 142 60 145
rect 68 142 70 145
rect 153 159 156 161
rect 167 152 169 155
rect 103 142 105 145
rect 113 142 115 145
rect 198 159 201 161
rect 212 152 214 155
rect 148 142 150 145
rect 158 142 160 145
rect 243 159 246 161
rect 257 152 259 155
rect 193 142 195 145
rect 203 142 205 145
rect 288 159 291 161
rect 302 152 304 155
rect 238 142 240 145
rect 248 142 250 145
rect 333 159 336 161
rect 347 152 349 155
rect 283 142 285 145
rect 293 142 295 145
rect 378 159 381 161
rect 392 152 394 155
rect 328 142 330 145
rect 338 142 340 145
rect 423 159 426 161
rect 437 152 439 155
rect 373 142 375 145
rect 383 142 385 145
rect 468 159 471 161
rect 482 152 484 155
rect 418 142 420 145
rect 428 142 430 145
rect 513 159 516 161
rect 527 152 529 155
rect 463 142 465 145
rect 473 142 475 145
rect 558 159 561 161
rect 572 152 574 155
rect 508 142 510 145
rect 518 142 520 145
rect 603 159 606 161
rect 617 152 619 155
rect 553 142 555 145
rect 563 142 565 145
rect 648 159 651 161
rect 662 152 664 155
rect 598 142 600 145
rect 608 142 610 145
rect 693 159 696 161
rect 707 152 709 155
rect 643 142 645 145
rect 653 142 655 145
rect 738 159 741 161
rect 752 152 754 155
rect 688 142 690 145
rect 698 142 700 145
rect 783 159 786 161
rect 797 152 799 155
rect 733 142 735 145
rect 743 142 745 145
rect 828 159 831 161
rect 842 152 844 155
rect 778 142 780 145
rect 788 142 790 145
rect 873 159 876 161
rect 887 152 889 155
rect 823 142 825 145
rect 833 142 835 145
rect 868 142 870 145
rect 878 142 880 145
rect 18 114 21 116
rect 32 107 34 110
rect 63 114 66 116
rect 77 107 79 110
rect 13 97 15 100
rect 23 97 25 100
rect 108 114 111 116
rect 122 107 124 110
rect 58 97 60 100
rect 68 97 70 100
rect 153 114 156 116
rect 167 107 169 110
rect 103 97 105 100
rect 113 97 115 100
rect 198 114 201 116
rect 212 107 214 110
rect 148 97 150 100
rect 158 97 160 100
rect 243 114 246 116
rect 257 107 259 110
rect 193 97 195 100
rect 203 97 205 100
rect 288 114 291 116
rect 302 107 304 110
rect 238 97 240 100
rect 248 97 250 100
rect 333 114 336 116
rect 347 107 349 110
rect 283 97 285 100
rect 293 97 295 100
rect 378 114 381 116
rect 392 107 394 110
rect 328 97 330 100
rect 338 97 340 100
rect 423 114 426 116
rect 437 107 439 110
rect 373 97 375 100
rect 383 97 385 100
rect 468 114 471 116
rect 482 107 484 110
rect 418 97 420 100
rect 428 97 430 100
rect 513 114 516 116
rect 527 107 529 110
rect 463 97 465 100
rect 473 97 475 100
rect 558 114 561 116
rect 572 107 574 110
rect 508 97 510 100
rect 518 97 520 100
rect 603 114 606 116
rect 617 107 619 110
rect 553 97 555 100
rect 563 97 565 100
rect 648 114 651 116
rect 662 107 664 110
rect 598 97 600 100
rect 608 97 610 100
rect 693 114 696 116
rect 707 107 709 110
rect 643 97 645 100
rect 653 97 655 100
rect 738 114 741 116
rect 752 107 754 110
rect 688 97 690 100
rect 698 97 700 100
rect 783 114 786 116
rect 797 107 799 110
rect 733 97 735 100
rect 743 97 745 100
rect 828 114 831 116
rect 842 107 844 110
rect 778 97 780 100
rect 788 97 790 100
rect 873 114 876 116
rect 887 107 889 110
rect 823 97 825 100
rect 833 97 835 100
rect 868 97 870 100
rect 878 97 880 100
rect 18 69 21 71
rect 32 62 34 65
rect 63 69 66 71
rect 77 62 79 65
rect 13 52 15 55
rect 23 52 25 55
rect 108 69 111 71
rect 122 62 124 65
rect 58 52 60 55
rect 68 52 70 55
rect 153 69 156 71
rect 167 62 169 65
rect 103 52 105 55
rect 113 52 115 55
rect 198 69 201 71
rect 212 62 214 65
rect 148 52 150 55
rect 158 52 160 55
rect 243 69 246 71
rect 257 62 259 65
rect 193 52 195 55
rect 203 52 205 55
rect 288 69 291 71
rect 302 62 304 65
rect 238 52 240 55
rect 248 52 250 55
rect 333 69 336 71
rect 347 62 349 65
rect 283 52 285 55
rect 293 52 295 55
rect 378 69 381 71
rect 392 62 394 65
rect 328 52 330 55
rect 338 52 340 55
rect 423 69 426 71
rect 437 62 439 65
rect 373 52 375 55
rect 383 52 385 55
rect 468 69 471 71
rect 482 62 484 65
rect 418 52 420 55
rect 428 52 430 55
rect 513 69 516 71
rect 527 62 529 65
rect 463 52 465 55
rect 473 52 475 55
rect 558 69 561 71
rect 572 62 574 65
rect 508 52 510 55
rect 518 52 520 55
rect 603 69 606 71
rect 617 62 619 65
rect 553 52 555 55
rect 563 52 565 55
rect 648 69 651 71
rect 662 62 664 65
rect 598 52 600 55
rect 608 52 610 55
rect 693 69 696 71
rect 707 62 709 65
rect 643 52 645 55
rect 653 52 655 55
rect 738 69 741 71
rect 752 62 754 65
rect 688 52 690 55
rect 698 52 700 55
rect 783 69 786 71
rect 797 62 799 65
rect 733 52 735 55
rect 743 52 745 55
rect 828 69 831 71
rect 842 62 844 65
rect 778 52 780 55
rect 788 52 790 55
rect 873 69 876 71
rect 887 62 889 65
rect 823 52 825 55
rect 833 52 835 55
rect 868 52 870 55
rect 878 52 880 55
rect 18 24 21 26
rect 32 17 34 20
rect 63 24 66 26
rect 77 17 79 20
rect 13 7 15 10
rect 23 7 25 10
rect 108 24 111 26
rect 122 17 124 20
rect 58 7 60 10
rect 68 7 70 10
rect 153 24 156 26
rect 167 17 169 20
rect 103 7 105 10
rect 113 7 115 10
rect 198 24 201 26
rect 212 17 214 20
rect 148 7 150 10
rect 158 7 160 10
rect 243 24 246 26
rect 257 17 259 20
rect 193 7 195 10
rect 203 7 205 10
rect 288 24 291 26
rect 302 17 304 20
rect 238 7 240 10
rect 248 7 250 10
rect 333 24 336 26
rect 347 17 349 20
rect 283 7 285 10
rect 293 7 295 10
rect 378 24 381 26
rect 392 17 394 20
rect 328 7 330 10
rect 338 7 340 10
rect 423 24 426 26
rect 437 17 439 20
rect 373 7 375 10
rect 383 7 385 10
rect 468 24 471 26
rect 482 17 484 20
rect 418 7 420 10
rect 428 7 430 10
rect 513 24 516 26
rect 527 17 529 20
rect 463 7 465 10
rect 473 7 475 10
rect 558 24 561 26
rect 572 17 574 20
rect 508 7 510 10
rect 518 7 520 10
rect 603 24 606 26
rect 617 17 619 20
rect 553 7 555 10
rect 563 7 565 10
rect 648 24 651 26
rect 662 17 664 20
rect 598 7 600 10
rect 608 7 610 10
rect 693 24 696 26
rect 707 17 709 20
rect 643 7 645 10
rect 653 7 655 10
rect 738 24 741 26
rect 752 17 754 20
rect 688 7 690 10
rect 698 7 700 10
rect 783 24 786 26
rect 797 17 799 20
rect 733 7 735 10
rect 743 7 745 10
rect 828 24 831 26
rect 842 17 844 20
rect 778 7 780 10
rect 788 7 790 10
rect 873 24 876 26
rect 887 17 889 20
rect 823 7 825 10
rect 833 7 835 10
rect 868 7 870 10
rect 878 7 880 10
rect -292 -169 -290 -163
rect -287 -169 -285 -163
rect -268 -165 -263 -163
rect -198 -157 -195 -155
rect -184 -164 -182 -161
rect -260 -176 -258 -170
rect -203 -174 -201 -171
rect -193 -174 -191 -171
<< ndiffusion >>
rect 3 883 45 900
rect 3 882 23 883
rect 3 870 13 882
rect 18 881 21 882
rect 18 878 21 879
rect 29 879 45 883
rect 35 875 45 879
rect 31 872 32 875
rect 34 872 45 875
rect 35 870 45 872
rect 48 883 90 900
rect 48 882 68 883
rect 48 870 58 882
rect 63 881 66 882
rect 63 878 66 879
rect 74 879 90 883
rect 80 875 90 879
rect 76 872 77 875
rect 79 872 90 875
rect 12 862 13 865
rect 15 862 23 865
rect 25 862 27 865
rect 39 864 45 870
rect 35 858 45 864
rect 80 870 90 872
rect 93 883 135 900
rect 93 882 113 883
rect 93 870 103 882
rect 108 881 111 882
rect 108 878 111 879
rect 119 879 135 883
rect 125 875 135 879
rect 121 872 122 875
rect 124 872 135 875
rect 57 862 58 865
rect 60 862 68 865
rect 70 862 72 865
rect 84 864 90 870
rect 80 858 90 864
rect 125 870 135 872
rect 138 883 180 900
rect 138 882 158 883
rect 138 870 148 882
rect 153 881 156 882
rect 153 878 156 879
rect 164 879 180 883
rect 170 875 180 879
rect 166 872 167 875
rect 169 872 180 875
rect 102 862 103 865
rect 105 862 113 865
rect 115 862 117 865
rect 129 864 135 870
rect 125 858 135 864
rect 170 870 180 872
rect 183 883 225 900
rect 183 882 203 883
rect 183 870 193 882
rect 198 881 201 882
rect 198 878 201 879
rect 209 879 225 883
rect 215 875 225 879
rect 211 872 212 875
rect 214 872 225 875
rect 147 862 148 865
rect 150 862 158 865
rect 160 862 162 865
rect 174 864 180 870
rect 170 858 180 864
rect 215 870 225 872
rect 228 883 270 900
rect 228 882 248 883
rect 228 870 238 882
rect 243 881 246 882
rect 243 878 246 879
rect 254 879 270 883
rect 260 875 270 879
rect 256 872 257 875
rect 259 872 270 875
rect 192 862 193 865
rect 195 862 203 865
rect 205 862 207 865
rect 219 864 225 870
rect 215 858 225 864
rect 260 870 270 872
rect 273 883 315 900
rect 273 882 293 883
rect 273 870 283 882
rect 288 881 291 882
rect 288 878 291 879
rect 299 879 315 883
rect 305 875 315 879
rect 301 872 302 875
rect 304 872 315 875
rect 237 862 238 865
rect 240 862 248 865
rect 250 862 252 865
rect 264 864 270 870
rect 260 858 270 864
rect 305 870 315 872
rect 318 883 360 900
rect 318 882 338 883
rect 318 870 328 882
rect 333 881 336 882
rect 333 878 336 879
rect 344 879 360 883
rect 350 875 360 879
rect 346 872 347 875
rect 349 872 360 875
rect 282 862 283 865
rect 285 862 293 865
rect 295 862 297 865
rect 309 864 315 870
rect 305 858 315 864
rect 350 870 360 872
rect 363 883 405 900
rect 363 882 383 883
rect 363 870 373 882
rect 378 881 381 882
rect 378 878 381 879
rect 389 879 405 883
rect 395 875 405 879
rect 391 872 392 875
rect 394 872 405 875
rect 327 862 328 865
rect 330 862 338 865
rect 340 862 342 865
rect 354 864 360 870
rect 350 858 360 864
rect 395 870 405 872
rect 408 883 450 900
rect 408 882 428 883
rect 408 870 418 882
rect 423 881 426 882
rect 423 878 426 879
rect 434 879 450 883
rect 440 875 450 879
rect 436 872 437 875
rect 439 872 450 875
rect 372 862 373 865
rect 375 862 383 865
rect 385 862 387 865
rect 399 864 405 870
rect 395 858 405 864
rect 440 870 450 872
rect 453 883 495 900
rect 453 882 473 883
rect 453 870 463 882
rect 468 881 471 882
rect 468 878 471 879
rect 479 879 495 883
rect 485 875 495 879
rect 481 872 482 875
rect 484 872 495 875
rect 417 862 418 865
rect 420 862 428 865
rect 430 862 432 865
rect 444 864 450 870
rect 440 858 450 864
rect 485 870 495 872
rect 498 883 540 900
rect 498 882 518 883
rect 498 870 508 882
rect 513 881 516 882
rect 513 878 516 879
rect 524 879 540 883
rect 530 875 540 879
rect 526 872 527 875
rect 529 872 540 875
rect 462 862 463 865
rect 465 862 473 865
rect 475 862 477 865
rect 489 864 495 870
rect 485 858 495 864
rect 530 870 540 872
rect 543 883 585 900
rect 543 882 563 883
rect 543 870 553 882
rect 558 881 561 882
rect 558 878 561 879
rect 569 879 585 883
rect 575 875 585 879
rect 571 872 572 875
rect 574 872 585 875
rect 507 862 508 865
rect 510 862 518 865
rect 520 862 522 865
rect 534 864 540 870
rect 530 858 540 864
rect 575 870 585 872
rect 588 883 630 900
rect 588 882 608 883
rect 588 870 598 882
rect 603 881 606 882
rect 603 878 606 879
rect 614 879 630 883
rect 620 875 630 879
rect 616 872 617 875
rect 619 872 630 875
rect 552 862 553 865
rect 555 862 563 865
rect 565 862 567 865
rect 579 864 585 870
rect 575 858 585 864
rect 620 870 630 872
rect 633 883 675 900
rect 633 882 653 883
rect 633 870 643 882
rect 648 881 651 882
rect 648 878 651 879
rect 659 879 675 883
rect 665 875 675 879
rect 661 872 662 875
rect 664 872 675 875
rect 597 862 598 865
rect 600 862 608 865
rect 610 862 612 865
rect 624 864 630 870
rect 620 858 630 864
rect 665 870 675 872
rect 678 883 720 900
rect 678 882 698 883
rect 678 870 688 882
rect 693 881 696 882
rect 693 878 696 879
rect 704 879 720 883
rect 710 875 720 879
rect 706 872 707 875
rect 709 872 720 875
rect 642 862 643 865
rect 645 862 653 865
rect 655 862 657 865
rect 669 864 675 870
rect 665 858 675 864
rect 710 870 720 872
rect 723 883 765 900
rect 723 882 743 883
rect 723 870 733 882
rect 738 881 741 882
rect 738 878 741 879
rect 749 879 765 883
rect 755 875 765 879
rect 751 872 752 875
rect 754 872 765 875
rect 687 862 688 865
rect 690 862 698 865
rect 700 862 702 865
rect 714 864 720 870
rect 710 858 720 864
rect 755 870 765 872
rect 768 883 810 900
rect 768 882 788 883
rect 768 870 778 882
rect 783 881 786 882
rect 783 878 786 879
rect 794 879 810 883
rect 800 875 810 879
rect 796 872 797 875
rect 799 872 810 875
rect 732 862 733 865
rect 735 862 743 865
rect 745 862 747 865
rect 759 864 765 870
rect 755 858 765 864
rect 800 870 810 872
rect 813 883 855 900
rect 813 882 833 883
rect 813 870 823 882
rect 828 881 831 882
rect 828 878 831 879
rect 839 879 855 883
rect 845 875 855 879
rect 841 872 842 875
rect 844 872 855 875
rect 777 862 778 865
rect 780 862 788 865
rect 790 862 792 865
rect 804 864 810 870
rect 800 858 810 864
rect 845 870 855 872
rect 858 883 900 900
rect 858 882 878 883
rect 858 870 868 882
rect 873 881 876 882
rect 873 878 876 879
rect 884 879 900 883
rect 890 875 900 879
rect 886 872 887 875
rect 889 872 900 875
rect 822 862 823 865
rect 825 862 833 865
rect 835 862 837 865
rect 849 864 855 870
rect 845 858 855 864
rect 890 870 900 872
rect 867 862 868 865
rect 870 862 878 865
rect 880 862 882 865
rect 894 864 900 870
rect 890 858 900 864
rect 3 838 45 855
rect 3 837 23 838
rect 3 825 13 837
rect 18 836 21 837
rect 18 833 21 834
rect 29 834 45 838
rect 35 830 45 834
rect 31 827 32 830
rect 34 827 45 830
rect 35 825 45 827
rect 48 838 90 855
rect 48 837 68 838
rect 48 825 58 837
rect 63 836 66 837
rect 63 833 66 834
rect 74 834 90 838
rect 80 830 90 834
rect 76 827 77 830
rect 79 827 90 830
rect 12 817 13 820
rect 15 817 23 820
rect 25 817 27 820
rect 39 819 45 825
rect 35 813 45 819
rect 80 825 90 827
rect 93 838 135 855
rect 93 837 113 838
rect 93 825 103 837
rect 108 836 111 837
rect 108 833 111 834
rect 119 834 135 838
rect 125 830 135 834
rect 121 827 122 830
rect 124 827 135 830
rect 57 817 58 820
rect 60 817 68 820
rect 70 817 72 820
rect 84 819 90 825
rect 80 813 90 819
rect 125 825 135 827
rect 138 838 180 855
rect 138 837 158 838
rect 138 825 148 837
rect 153 836 156 837
rect 153 833 156 834
rect 164 834 180 838
rect 170 830 180 834
rect 166 827 167 830
rect 169 827 180 830
rect 102 817 103 820
rect 105 817 113 820
rect 115 817 117 820
rect 129 819 135 825
rect 125 813 135 819
rect 170 825 180 827
rect 183 838 225 855
rect 183 837 203 838
rect 183 825 193 837
rect 198 836 201 837
rect 198 833 201 834
rect 209 834 225 838
rect 215 830 225 834
rect 211 827 212 830
rect 214 827 225 830
rect 147 817 148 820
rect 150 817 158 820
rect 160 817 162 820
rect 174 819 180 825
rect 170 813 180 819
rect 215 825 225 827
rect 228 838 270 855
rect 228 837 248 838
rect 228 825 238 837
rect 243 836 246 837
rect 243 833 246 834
rect 254 834 270 838
rect 260 830 270 834
rect 256 827 257 830
rect 259 827 270 830
rect 192 817 193 820
rect 195 817 203 820
rect 205 817 207 820
rect 219 819 225 825
rect 215 813 225 819
rect 260 825 270 827
rect 273 838 315 855
rect 273 837 293 838
rect 273 825 283 837
rect 288 836 291 837
rect 288 833 291 834
rect 299 834 315 838
rect 305 830 315 834
rect 301 827 302 830
rect 304 827 315 830
rect 237 817 238 820
rect 240 817 248 820
rect 250 817 252 820
rect 264 819 270 825
rect 260 813 270 819
rect 305 825 315 827
rect 318 838 360 855
rect 318 837 338 838
rect 318 825 328 837
rect 333 836 336 837
rect 333 833 336 834
rect 344 834 360 838
rect 350 830 360 834
rect 346 827 347 830
rect 349 827 360 830
rect 282 817 283 820
rect 285 817 293 820
rect 295 817 297 820
rect 309 819 315 825
rect 305 813 315 819
rect 350 825 360 827
rect 363 838 405 855
rect 363 837 383 838
rect 363 825 373 837
rect 378 836 381 837
rect 378 833 381 834
rect 389 834 405 838
rect 395 830 405 834
rect 391 827 392 830
rect 394 827 405 830
rect 327 817 328 820
rect 330 817 338 820
rect 340 817 342 820
rect 354 819 360 825
rect 350 813 360 819
rect 395 825 405 827
rect 408 838 450 855
rect 408 837 428 838
rect 408 825 418 837
rect 423 836 426 837
rect 423 833 426 834
rect 434 834 450 838
rect 440 830 450 834
rect 436 827 437 830
rect 439 827 450 830
rect 372 817 373 820
rect 375 817 383 820
rect 385 817 387 820
rect 399 819 405 825
rect 395 813 405 819
rect 440 825 450 827
rect 453 838 495 855
rect 453 837 473 838
rect 453 825 463 837
rect 468 836 471 837
rect 468 833 471 834
rect 479 834 495 838
rect 485 830 495 834
rect 481 827 482 830
rect 484 827 495 830
rect 417 817 418 820
rect 420 817 428 820
rect 430 817 432 820
rect 444 819 450 825
rect 440 813 450 819
rect 485 825 495 827
rect 498 838 540 855
rect 498 837 518 838
rect 498 825 508 837
rect 513 836 516 837
rect 513 833 516 834
rect 524 834 540 838
rect 530 830 540 834
rect 526 827 527 830
rect 529 827 540 830
rect 462 817 463 820
rect 465 817 473 820
rect 475 817 477 820
rect 489 819 495 825
rect 485 813 495 819
rect 530 825 540 827
rect 543 838 585 855
rect 543 837 563 838
rect 543 825 553 837
rect 558 836 561 837
rect 558 833 561 834
rect 569 834 585 838
rect 575 830 585 834
rect 571 827 572 830
rect 574 827 585 830
rect 507 817 508 820
rect 510 817 518 820
rect 520 817 522 820
rect 534 819 540 825
rect 530 813 540 819
rect 575 825 585 827
rect 588 838 630 855
rect 588 837 608 838
rect 588 825 598 837
rect 603 836 606 837
rect 603 833 606 834
rect 614 834 630 838
rect 620 830 630 834
rect 616 827 617 830
rect 619 827 630 830
rect 552 817 553 820
rect 555 817 563 820
rect 565 817 567 820
rect 579 819 585 825
rect 575 813 585 819
rect 620 825 630 827
rect 633 838 675 855
rect 633 837 653 838
rect 633 825 643 837
rect 648 836 651 837
rect 648 833 651 834
rect 659 834 675 838
rect 665 830 675 834
rect 661 827 662 830
rect 664 827 675 830
rect 597 817 598 820
rect 600 817 608 820
rect 610 817 612 820
rect 624 819 630 825
rect 620 813 630 819
rect 665 825 675 827
rect 678 838 720 855
rect 678 837 698 838
rect 678 825 688 837
rect 693 836 696 837
rect 693 833 696 834
rect 704 834 720 838
rect 710 830 720 834
rect 706 827 707 830
rect 709 827 720 830
rect 642 817 643 820
rect 645 817 653 820
rect 655 817 657 820
rect 669 819 675 825
rect 665 813 675 819
rect 710 825 720 827
rect 723 838 765 855
rect 723 837 743 838
rect 723 825 733 837
rect 738 836 741 837
rect 738 833 741 834
rect 749 834 765 838
rect 755 830 765 834
rect 751 827 752 830
rect 754 827 765 830
rect 687 817 688 820
rect 690 817 698 820
rect 700 817 702 820
rect 714 819 720 825
rect 710 813 720 819
rect 755 825 765 827
rect 768 838 810 855
rect 768 837 788 838
rect 768 825 778 837
rect 783 836 786 837
rect 783 833 786 834
rect 794 834 810 838
rect 800 830 810 834
rect 796 827 797 830
rect 799 827 810 830
rect 732 817 733 820
rect 735 817 743 820
rect 745 817 747 820
rect 759 819 765 825
rect 755 813 765 819
rect 800 825 810 827
rect 813 838 855 855
rect 813 837 833 838
rect 813 825 823 837
rect 828 836 831 837
rect 828 833 831 834
rect 839 834 855 838
rect 845 830 855 834
rect 841 827 842 830
rect 844 827 855 830
rect 777 817 778 820
rect 780 817 788 820
rect 790 817 792 820
rect 804 819 810 825
rect 800 813 810 819
rect 845 825 855 827
rect 858 838 900 855
rect 858 837 878 838
rect 858 825 868 837
rect 873 836 876 837
rect 873 833 876 834
rect 884 834 900 838
rect 890 830 900 834
rect 886 827 887 830
rect 889 827 900 830
rect 822 817 823 820
rect 825 817 833 820
rect 835 817 837 820
rect 849 819 855 825
rect 845 813 855 819
rect 890 825 900 827
rect 867 817 868 820
rect 870 817 878 820
rect 880 817 882 820
rect 894 819 900 825
rect 890 813 900 819
rect 3 793 45 810
rect 3 792 23 793
rect 3 780 13 792
rect 18 791 21 792
rect 18 788 21 789
rect 29 789 45 793
rect 35 785 45 789
rect 31 782 32 785
rect 34 782 45 785
rect 35 780 45 782
rect 48 793 90 810
rect 48 792 68 793
rect 48 780 58 792
rect 63 791 66 792
rect 63 788 66 789
rect 74 789 90 793
rect 80 785 90 789
rect 76 782 77 785
rect 79 782 90 785
rect 12 772 13 775
rect 15 772 23 775
rect 25 772 27 775
rect 39 774 45 780
rect 35 768 45 774
rect 80 780 90 782
rect 93 793 135 810
rect 93 792 113 793
rect 93 780 103 792
rect 108 791 111 792
rect 108 788 111 789
rect 119 789 135 793
rect 125 785 135 789
rect 121 782 122 785
rect 124 782 135 785
rect 57 772 58 775
rect 60 772 68 775
rect 70 772 72 775
rect 84 774 90 780
rect 80 768 90 774
rect 125 780 135 782
rect 138 793 180 810
rect 138 792 158 793
rect 138 780 148 792
rect 153 791 156 792
rect 153 788 156 789
rect 164 789 180 793
rect 170 785 180 789
rect 166 782 167 785
rect 169 782 180 785
rect 102 772 103 775
rect 105 772 113 775
rect 115 772 117 775
rect 129 774 135 780
rect 125 768 135 774
rect 170 780 180 782
rect 183 793 225 810
rect 183 792 203 793
rect 183 780 193 792
rect 198 791 201 792
rect 198 788 201 789
rect 209 789 225 793
rect 215 785 225 789
rect 211 782 212 785
rect 214 782 225 785
rect 147 772 148 775
rect 150 772 158 775
rect 160 772 162 775
rect 174 774 180 780
rect 170 768 180 774
rect 215 780 225 782
rect 228 793 270 810
rect 228 792 248 793
rect 228 780 238 792
rect 243 791 246 792
rect 243 788 246 789
rect 254 789 270 793
rect 260 785 270 789
rect 256 782 257 785
rect 259 782 270 785
rect 192 772 193 775
rect 195 772 203 775
rect 205 772 207 775
rect 219 774 225 780
rect 215 768 225 774
rect 260 780 270 782
rect 273 793 315 810
rect 273 792 293 793
rect 273 780 283 792
rect 288 791 291 792
rect 288 788 291 789
rect 299 789 315 793
rect 305 785 315 789
rect 301 782 302 785
rect 304 782 315 785
rect 237 772 238 775
rect 240 772 248 775
rect 250 772 252 775
rect 264 774 270 780
rect 260 768 270 774
rect 305 780 315 782
rect 318 793 360 810
rect 318 792 338 793
rect 318 780 328 792
rect 333 791 336 792
rect 333 788 336 789
rect 344 789 360 793
rect 350 785 360 789
rect 346 782 347 785
rect 349 782 360 785
rect 282 772 283 775
rect 285 772 293 775
rect 295 772 297 775
rect 309 774 315 780
rect 305 768 315 774
rect 350 780 360 782
rect 363 793 405 810
rect 363 792 383 793
rect 363 780 373 792
rect 378 791 381 792
rect 378 788 381 789
rect 389 789 405 793
rect 395 785 405 789
rect 391 782 392 785
rect 394 782 405 785
rect 327 772 328 775
rect 330 772 338 775
rect 340 772 342 775
rect 354 774 360 780
rect 350 768 360 774
rect 395 780 405 782
rect 408 793 450 810
rect 408 792 428 793
rect 408 780 418 792
rect 423 791 426 792
rect 423 788 426 789
rect 434 789 450 793
rect 440 785 450 789
rect 436 782 437 785
rect 439 782 450 785
rect 372 772 373 775
rect 375 772 383 775
rect 385 772 387 775
rect 399 774 405 780
rect 395 768 405 774
rect 440 780 450 782
rect 453 793 495 810
rect 453 792 473 793
rect 453 780 463 792
rect 468 791 471 792
rect 468 788 471 789
rect 479 789 495 793
rect 485 785 495 789
rect 481 782 482 785
rect 484 782 495 785
rect 417 772 418 775
rect 420 772 428 775
rect 430 772 432 775
rect 444 774 450 780
rect 440 768 450 774
rect 485 780 495 782
rect 498 793 540 810
rect 498 792 518 793
rect 498 780 508 792
rect 513 791 516 792
rect 513 788 516 789
rect 524 789 540 793
rect 530 785 540 789
rect 526 782 527 785
rect 529 782 540 785
rect 462 772 463 775
rect 465 772 473 775
rect 475 772 477 775
rect 489 774 495 780
rect 485 768 495 774
rect 530 780 540 782
rect 543 793 585 810
rect 543 792 563 793
rect 543 780 553 792
rect 558 791 561 792
rect 558 788 561 789
rect 569 789 585 793
rect 575 785 585 789
rect 571 782 572 785
rect 574 782 585 785
rect 507 772 508 775
rect 510 772 518 775
rect 520 772 522 775
rect 534 774 540 780
rect 530 768 540 774
rect 575 780 585 782
rect 588 793 630 810
rect 588 792 608 793
rect 588 780 598 792
rect 603 791 606 792
rect 603 788 606 789
rect 614 789 630 793
rect 620 785 630 789
rect 616 782 617 785
rect 619 782 630 785
rect 552 772 553 775
rect 555 772 563 775
rect 565 772 567 775
rect 579 774 585 780
rect 575 768 585 774
rect 620 780 630 782
rect 633 793 675 810
rect 633 792 653 793
rect 633 780 643 792
rect 648 791 651 792
rect 648 788 651 789
rect 659 789 675 793
rect 665 785 675 789
rect 661 782 662 785
rect 664 782 675 785
rect 597 772 598 775
rect 600 772 608 775
rect 610 772 612 775
rect 624 774 630 780
rect 620 768 630 774
rect 665 780 675 782
rect 678 793 720 810
rect 678 792 698 793
rect 678 780 688 792
rect 693 791 696 792
rect 693 788 696 789
rect 704 789 720 793
rect 710 785 720 789
rect 706 782 707 785
rect 709 782 720 785
rect 642 772 643 775
rect 645 772 653 775
rect 655 772 657 775
rect 669 774 675 780
rect 665 768 675 774
rect 710 780 720 782
rect 723 793 765 810
rect 723 792 743 793
rect 723 780 733 792
rect 738 791 741 792
rect 738 788 741 789
rect 749 789 765 793
rect 755 785 765 789
rect 751 782 752 785
rect 754 782 765 785
rect 687 772 688 775
rect 690 772 698 775
rect 700 772 702 775
rect 714 774 720 780
rect 710 768 720 774
rect 755 780 765 782
rect 768 793 810 810
rect 768 792 788 793
rect 768 780 778 792
rect 783 791 786 792
rect 783 788 786 789
rect 794 789 810 793
rect 800 785 810 789
rect 796 782 797 785
rect 799 782 810 785
rect 732 772 733 775
rect 735 772 743 775
rect 745 772 747 775
rect 759 774 765 780
rect 755 768 765 774
rect 800 780 810 782
rect 813 793 855 810
rect 813 792 833 793
rect 813 780 823 792
rect 828 791 831 792
rect 828 788 831 789
rect 839 789 855 793
rect 845 785 855 789
rect 841 782 842 785
rect 844 782 855 785
rect 777 772 778 775
rect 780 772 788 775
rect 790 772 792 775
rect 804 774 810 780
rect 800 768 810 774
rect 845 780 855 782
rect 858 793 900 810
rect 858 792 878 793
rect 858 780 868 792
rect 873 791 876 792
rect 873 788 876 789
rect 884 789 900 793
rect 890 785 900 789
rect 886 782 887 785
rect 889 782 900 785
rect 822 772 823 775
rect 825 772 833 775
rect 835 772 837 775
rect 849 774 855 780
rect 845 768 855 774
rect 890 780 900 782
rect 867 772 868 775
rect 870 772 878 775
rect 880 772 882 775
rect 894 774 900 780
rect 890 768 900 774
rect 3 748 45 765
rect 3 747 23 748
rect 3 735 13 747
rect 18 746 21 747
rect 18 743 21 744
rect 29 744 45 748
rect 35 740 45 744
rect 31 737 32 740
rect 34 737 45 740
rect 35 735 45 737
rect 48 748 90 765
rect 48 747 68 748
rect 48 735 58 747
rect 63 746 66 747
rect 63 743 66 744
rect 74 744 90 748
rect 80 740 90 744
rect 76 737 77 740
rect 79 737 90 740
rect 12 727 13 730
rect 15 727 23 730
rect 25 727 27 730
rect 39 729 45 735
rect 35 723 45 729
rect 80 735 90 737
rect 93 748 135 765
rect 93 747 113 748
rect 93 735 103 747
rect 108 746 111 747
rect 108 743 111 744
rect 119 744 135 748
rect 125 740 135 744
rect 121 737 122 740
rect 124 737 135 740
rect 57 727 58 730
rect 60 727 68 730
rect 70 727 72 730
rect 84 729 90 735
rect 80 723 90 729
rect 125 735 135 737
rect 138 748 180 765
rect 138 747 158 748
rect 138 735 148 747
rect 153 746 156 747
rect 153 743 156 744
rect 164 744 180 748
rect 170 740 180 744
rect 166 737 167 740
rect 169 737 180 740
rect 102 727 103 730
rect 105 727 113 730
rect 115 727 117 730
rect 129 729 135 735
rect 125 723 135 729
rect 170 735 180 737
rect 183 748 225 765
rect 183 747 203 748
rect 183 735 193 747
rect 198 746 201 747
rect 198 743 201 744
rect 209 744 225 748
rect 215 740 225 744
rect 211 737 212 740
rect 214 737 225 740
rect 147 727 148 730
rect 150 727 158 730
rect 160 727 162 730
rect 174 729 180 735
rect 170 723 180 729
rect 215 735 225 737
rect 228 748 270 765
rect 228 747 248 748
rect 228 735 238 747
rect 243 746 246 747
rect 243 743 246 744
rect 254 744 270 748
rect 260 740 270 744
rect 256 737 257 740
rect 259 737 270 740
rect 192 727 193 730
rect 195 727 203 730
rect 205 727 207 730
rect 219 729 225 735
rect 215 723 225 729
rect 260 735 270 737
rect 273 748 315 765
rect 273 747 293 748
rect 273 735 283 747
rect 288 746 291 747
rect 288 743 291 744
rect 299 744 315 748
rect 305 740 315 744
rect 301 737 302 740
rect 304 737 315 740
rect 237 727 238 730
rect 240 727 248 730
rect 250 727 252 730
rect 264 729 270 735
rect 260 723 270 729
rect 305 735 315 737
rect 318 748 360 765
rect 318 747 338 748
rect 318 735 328 747
rect 333 746 336 747
rect 333 743 336 744
rect 344 744 360 748
rect 350 740 360 744
rect 346 737 347 740
rect 349 737 360 740
rect 282 727 283 730
rect 285 727 293 730
rect 295 727 297 730
rect 309 729 315 735
rect 305 723 315 729
rect 350 735 360 737
rect 363 748 405 765
rect 363 747 383 748
rect 363 735 373 747
rect 378 746 381 747
rect 378 743 381 744
rect 389 744 405 748
rect 395 740 405 744
rect 391 737 392 740
rect 394 737 405 740
rect 327 727 328 730
rect 330 727 338 730
rect 340 727 342 730
rect 354 729 360 735
rect 350 723 360 729
rect 395 735 405 737
rect 408 748 450 765
rect 408 747 428 748
rect 408 735 418 747
rect 423 746 426 747
rect 423 743 426 744
rect 434 744 450 748
rect 440 740 450 744
rect 436 737 437 740
rect 439 737 450 740
rect 372 727 373 730
rect 375 727 383 730
rect 385 727 387 730
rect 399 729 405 735
rect 395 723 405 729
rect 440 735 450 737
rect 453 748 495 765
rect 453 747 473 748
rect 453 735 463 747
rect 468 746 471 747
rect 468 743 471 744
rect 479 744 495 748
rect 485 740 495 744
rect 481 737 482 740
rect 484 737 495 740
rect 417 727 418 730
rect 420 727 428 730
rect 430 727 432 730
rect 444 729 450 735
rect 440 723 450 729
rect 485 735 495 737
rect 498 748 540 765
rect 498 747 518 748
rect 498 735 508 747
rect 513 746 516 747
rect 513 743 516 744
rect 524 744 540 748
rect 530 740 540 744
rect 526 737 527 740
rect 529 737 540 740
rect 462 727 463 730
rect 465 727 473 730
rect 475 727 477 730
rect 489 729 495 735
rect 485 723 495 729
rect 530 735 540 737
rect 543 748 585 765
rect 543 747 563 748
rect 543 735 553 747
rect 558 746 561 747
rect 558 743 561 744
rect 569 744 585 748
rect 575 740 585 744
rect 571 737 572 740
rect 574 737 585 740
rect 507 727 508 730
rect 510 727 518 730
rect 520 727 522 730
rect 534 729 540 735
rect 530 723 540 729
rect 575 735 585 737
rect 588 748 630 765
rect 588 747 608 748
rect 588 735 598 747
rect 603 746 606 747
rect 603 743 606 744
rect 614 744 630 748
rect 620 740 630 744
rect 616 737 617 740
rect 619 737 630 740
rect 552 727 553 730
rect 555 727 563 730
rect 565 727 567 730
rect 579 729 585 735
rect 575 723 585 729
rect 620 735 630 737
rect 633 748 675 765
rect 633 747 653 748
rect 633 735 643 747
rect 648 746 651 747
rect 648 743 651 744
rect 659 744 675 748
rect 665 740 675 744
rect 661 737 662 740
rect 664 737 675 740
rect 597 727 598 730
rect 600 727 608 730
rect 610 727 612 730
rect 624 729 630 735
rect 620 723 630 729
rect 665 735 675 737
rect 678 748 720 765
rect 678 747 698 748
rect 678 735 688 747
rect 693 746 696 747
rect 693 743 696 744
rect 704 744 720 748
rect 710 740 720 744
rect 706 737 707 740
rect 709 737 720 740
rect 642 727 643 730
rect 645 727 653 730
rect 655 727 657 730
rect 669 729 675 735
rect 665 723 675 729
rect 710 735 720 737
rect 723 748 765 765
rect 723 747 743 748
rect 723 735 733 747
rect 738 746 741 747
rect 738 743 741 744
rect 749 744 765 748
rect 755 740 765 744
rect 751 737 752 740
rect 754 737 765 740
rect 687 727 688 730
rect 690 727 698 730
rect 700 727 702 730
rect 714 729 720 735
rect 710 723 720 729
rect 755 735 765 737
rect 768 748 810 765
rect 768 747 788 748
rect 768 735 778 747
rect 783 746 786 747
rect 783 743 786 744
rect 794 744 810 748
rect 800 740 810 744
rect 796 737 797 740
rect 799 737 810 740
rect 732 727 733 730
rect 735 727 743 730
rect 745 727 747 730
rect 759 729 765 735
rect 755 723 765 729
rect 800 735 810 737
rect 813 748 855 765
rect 813 747 833 748
rect 813 735 823 747
rect 828 746 831 747
rect 828 743 831 744
rect 839 744 855 748
rect 845 740 855 744
rect 841 737 842 740
rect 844 737 855 740
rect 777 727 778 730
rect 780 727 788 730
rect 790 727 792 730
rect 804 729 810 735
rect 800 723 810 729
rect 845 735 855 737
rect 858 748 900 765
rect 858 747 878 748
rect 858 735 868 747
rect 873 746 876 747
rect 873 743 876 744
rect 884 744 900 748
rect 890 740 900 744
rect 886 737 887 740
rect 889 737 900 740
rect 822 727 823 730
rect 825 727 833 730
rect 835 727 837 730
rect 849 729 855 735
rect 845 723 855 729
rect 890 735 900 737
rect 867 727 868 730
rect 870 727 878 730
rect 880 727 882 730
rect 894 729 900 735
rect 890 723 900 729
rect 3 703 45 720
rect 3 702 23 703
rect 3 690 13 702
rect 18 701 21 702
rect 18 698 21 699
rect 29 699 45 703
rect 35 695 45 699
rect 31 692 32 695
rect 34 692 45 695
rect 35 690 45 692
rect 48 703 90 720
rect 48 702 68 703
rect 48 690 58 702
rect 63 701 66 702
rect 63 698 66 699
rect 74 699 90 703
rect 80 695 90 699
rect 76 692 77 695
rect 79 692 90 695
rect 12 682 13 685
rect 15 682 23 685
rect 25 682 27 685
rect 39 684 45 690
rect 35 678 45 684
rect 80 690 90 692
rect 93 703 135 720
rect 93 702 113 703
rect 93 690 103 702
rect 108 701 111 702
rect 108 698 111 699
rect 119 699 135 703
rect 125 695 135 699
rect 121 692 122 695
rect 124 692 135 695
rect 57 682 58 685
rect 60 682 68 685
rect 70 682 72 685
rect 84 684 90 690
rect 80 678 90 684
rect 125 690 135 692
rect 138 703 180 720
rect 138 702 158 703
rect 138 690 148 702
rect 153 701 156 702
rect 153 698 156 699
rect 164 699 180 703
rect 170 695 180 699
rect 166 692 167 695
rect 169 692 180 695
rect 102 682 103 685
rect 105 682 113 685
rect 115 682 117 685
rect 129 684 135 690
rect 125 678 135 684
rect 170 690 180 692
rect 183 703 225 720
rect 183 702 203 703
rect 183 690 193 702
rect 198 701 201 702
rect 198 698 201 699
rect 209 699 225 703
rect 215 695 225 699
rect 211 692 212 695
rect 214 692 225 695
rect 147 682 148 685
rect 150 682 158 685
rect 160 682 162 685
rect 174 684 180 690
rect 170 678 180 684
rect 215 690 225 692
rect 228 703 270 720
rect 228 702 248 703
rect 228 690 238 702
rect 243 701 246 702
rect 243 698 246 699
rect 254 699 270 703
rect 260 695 270 699
rect 256 692 257 695
rect 259 692 270 695
rect 192 682 193 685
rect 195 682 203 685
rect 205 682 207 685
rect 219 684 225 690
rect 215 678 225 684
rect 260 690 270 692
rect 273 703 315 720
rect 273 702 293 703
rect 273 690 283 702
rect 288 701 291 702
rect 288 698 291 699
rect 299 699 315 703
rect 305 695 315 699
rect 301 692 302 695
rect 304 692 315 695
rect 237 682 238 685
rect 240 682 248 685
rect 250 682 252 685
rect 264 684 270 690
rect 260 678 270 684
rect 305 690 315 692
rect 318 703 360 720
rect 318 702 338 703
rect 318 690 328 702
rect 333 701 336 702
rect 333 698 336 699
rect 344 699 360 703
rect 350 695 360 699
rect 346 692 347 695
rect 349 692 360 695
rect 282 682 283 685
rect 285 682 293 685
rect 295 682 297 685
rect 309 684 315 690
rect 305 678 315 684
rect 350 690 360 692
rect 363 703 405 720
rect 363 702 383 703
rect 363 690 373 702
rect 378 701 381 702
rect 378 698 381 699
rect 389 699 405 703
rect 395 695 405 699
rect 391 692 392 695
rect 394 692 405 695
rect 327 682 328 685
rect 330 682 338 685
rect 340 682 342 685
rect 354 684 360 690
rect 350 678 360 684
rect 395 690 405 692
rect 408 703 450 720
rect 408 702 428 703
rect 408 690 418 702
rect 423 701 426 702
rect 423 698 426 699
rect 434 699 450 703
rect 440 695 450 699
rect 436 692 437 695
rect 439 692 450 695
rect 372 682 373 685
rect 375 682 383 685
rect 385 682 387 685
rect 399 684 405 690
rect 395 678 405 684
rect 440 690 450 692
rect 453 703 495 720
rect 453 702 473 703
rect 453 690 463 702
rect 468 701 471 702
rect 468 698 471 699
rect 479 699 495 703
rect 485 695 495 699
rect 481 692 482 695
rect 484 692 495 695
rect 417 682 418 685
rect 420 682 428 685
rect 430 682 432 685
rect 444 684 450 690
rect 440 678 450 684
rect 485 690 495 692
rect 498 703 540 720
rect 498 702 518 703
rect 498 690 508 702
rect 513 701 516 702
rect 513 698 516 699
rect 524 699 540 703
rect 530 695 540 699
rect 526 692 527 695
rect 529 692 540 695
rect 462 682 463 685
rect 465 682 473 685
rect 475 682 477 685
rect 489 684 495 690
rect 485 678 495 684
rect 530 690 540 692
rect 543 703 585 720
rect 543 702 563 703
rect 543 690 553 702
rect 558 701 561 702
rect 558 698 561 699
rect 569 699 585 703
rect 575 695 585 699
rect 571 692 572 695
rect 574 692 585 695
rect 507 682 508 685
rect 510 682 518 685
rect 520 682 522 685
rect 534 684 540 690
rect 530 678 540 684
rect 575 690 585 692
rect 588 703 630 720
rect 588 702 608 703
rect 588 690 598 702
rect 603 701 606 702
rect 603 698 606 699
rect 614 699 630 703
rect 620 695 630 699
rect 616 692 617 695
rect 619 692 630 695
rect 552 682 553 685
rect 555 682 563 685
rect 565 682 567 685
rect 579 684 585 690
rect 575 678 585 684
rect 620 690 630 692
rect 633 703 675 720
rect 633 702 653 703
rect 633 690 643 702
rect 648 701 651 702
rect 648 698 651 699
rect 659 699 675 703
rect 665 695 675 699
rect 661 692 662 695
rect 664 692 675 695
rect 597 682 598 685
rect 600 682 608 685
rect 610 682 612 685
rect 624 684 630 690
rect 620 678 630 684
rect 665 690 675 692
rect 678 703 720 720
rect 678 702 698 703
rect 678 690 688 702
rect 693 701 696 702
rect 693 698 696 699
rect 704 699 720 703
rect 710 695 720 699
rect 706 692 707 695
rect 709 692 720 695
rect 642 682 643 685
rect 645 682 653 685
rect 655 682 657 685
rect 669 684 675 690
rect 665 678 675 684
rect 710 690 720 692
rect 723 703 765 720
rect 723 702 743 703
rect 723 690 733 702
rect 738 701 741 702
rect 738 698 741 699
rect 749 699 765 703
rect 755 695 765 699
rect 751 692 752 695
rect 754 692 765 695
rect 687 682 688 685
rect 690 682 698 685
rect 700 682 702 685
rect 714 684 720 690
rect 710 678 720 684
rect 755 690 765 692
rect 768 703 810 720
rect 768 702 788 703
rect 768 690 778 702
rect 783 701 786 702
rect 783 698 786 699
rect 794 699 810 703
rect 800 695 810 699
rect 796 692 797 695
rect 799 692 810 695
rect 732 682 733 685
rect 735 682 743 685
rect 745 682 747 685
rect 759 684 765 690
rect 755 678 765 684
rect 800 690 810 692
rect 813 703 855 720
rect 813 702 833 703
rect 813 690 823 702
rect 828 701 831 702
rect 828 698 831 699
rect 839 699 855 703
rect 845 695 855 699
rect 841 692 842 695
rect 844 692 855 695
rect 777 682 778 685
rect 780 682 788 685
rect 790 682 792 685
rect 804 684 810 690
rect 800 678 810 684
rect 845 690 855 692
rect 858 703 900 720
rect 858 702 878 703
rect 858 690 868 702
rect 873 701 876 702
rect 873 698 876 699
rect 884 699 900 703
rect 890 695 900 699
rect 886 692 887 695
rect 889 692 900 695
rect 822 682 823 685
rect 825 682 833 685
rect 835 682 837 685
rect 849 684 855 690
rect 845 678 855 684
rect 890 690 900 692
rect 867 682 868 685
rect 870 682 878 685
rect 880 682 882 685
rect 894 684 900 690
rect 890 678 900 684
rect 3 658 45 675
rect 3 657 23 658
rect 3 645 13 657
rect 18 656 21 657
rect 18 653 21 654
rect 29 654 45 658
rect 35 650 45 654
rect 31 647 32 650
rect 34 647 45 650
rect 35 645 45 647
rect 48 658 90 675
rect 48 657 68 658
rect 48 645 58 657
rect 63 656 66 657
rect 63 653 66 654
rect 74 654 90 658
rect 80 650 90 654
rect 76 647 77 650
rect 79 647 90 650
rect 12 637 13 640
rect 15 637 23 640
rect 25 637 27 640
rect 39 639 45 645
rect 35 633 45 639
rect 80 645 90 647
rect 93 658 135 675
rect 93 657 113 658
rect 93 645 103 657
rect 108 656 111 657
rect 108 653 111 654
rect 119 654 135 658
rect 125 650 135 654
rect 121 647 122 650
rect 124 647 135 650
rect 57 637 58 640
rect 60 637 68 640
rect 70 637 72 640
rect 84 639 90 645
rect 80 633 90 639
rect 125 645 135 647
rect 138 658 180 675
rect 138 657 158 658
rect 138 645 148 657
rect 153 656 156 657
rect 153 653 156 654
rect 164 654 180 658
rect 170 650 180 654
rect 166 647 167 650
rect 169 647 180 650
rect 102 637 103 640
rect 105 637 113 640
rect 115 637 117 640
rect 129 639 135 645
rect 125 633 135 639
rect 170 645 180 647
rect 183 658 225 675
rect 183 657 203 658
rect 183 645 193 657
rect 198 656 201 657
rect 198 653 201 654
rect 209 654 225 658
rect 215 650 225 654
rect 211 647 212 650
rect 214 647 225 650
rect 147 637 148 640
rect 150 637 158 640
rect 160 637 162 640
rect 174 639 180 645
rect 170 633 180 639
rect 215 645 225 647
rect 228 658 270 675
rect 228 657 248 658
rect 228 645 238 657
rect 243 656 246 657
rect 243 653 246 654
rect 254 654 270 658
rect 260 650 270 654
rect 256 647 257 650
rect 259 647 270 650
rect 192 637 193 640
rect 195 637 203 640
rect 205 637 207 640
rect 219 639 225 645
rect 215 633 225 639
rect 260 645 270 647
rect 273 658 315 675
rect 273 657 293 658
rect 273 645 283 657
rect 288 656 291 657
rect 288 653 291 654
rect 299 654 315 658
rect 305 650 315 654
rect 301 647 302 650
rect 304 647 315 650
rect 237 637 238 640
rect 240 637 248 640
rect 250 637 252 640
rect 264 639 270 645
rect 260 633 270 639
rect 305 645 315 647
rect 318 658 360 675
rect 318 657 338 658
rect 318 645 328 657
rect 333 656 336 657
rect 333 653 336 654
rect 344 654 360 658
rect 350 650 360 654
rect 346 647 347 650
rect 349 647 360 650
rect 282 637 283 640
rect 285 637 293 640
rect 295 637 297 640
rect 309 639 315 645
rect 305 633 315 639
rect 350 645 360 647
rect 363 658 405 675
rect 363 657 383 658
rect 363 645 373 657
rect 378 656 381 657
rect 378 653 381 654
rect 389 654 405 658
rect 395 650 405 654
rect 391 647 392 650
rect 394 647 405 650
rect 327 637 328 640
rect 330 637 338 640
rect 340 637 342 640
rect 354 639 360 645
rect 350 633 360 639
rect 395 645 405 647
rect 408 658 450 675
rect 408 657 428 658
rect 408 645 418 657
rect 423 656 426 657
rect 423 653 426 654
rect 434 654 450 658
rect 440 650 450 654
rect 436 647 437 650
rect 439 647 450 650
rect 372 637 373 640
rect 375 637 383 640
rect 385 637 387 640
rect 399 639 405 645
rect 395 633 405 639
rect 440 645 450 647
rect 453 658 495 675
rect 453 657 473 658
rect 453 645 463 657
rect 468 656 471 657
rect 468 653 471 654
rect 479 654 495 658
rect 485 650 495 654
rect 481 647 482 650
rect 484 647 495 650
rect 417 637 418 640
rect 420 637 428 640
rect 430 637 432 640
rect 444 639 450 645
rect 440 633 450 639
rect 485 645 495 647
rect 498 658 540 675
rect 498 657 518 658
rect 498 645 508 657
rect 513 656 516 657
rect 513 653 516 654
rect 524 654 540 658
rect 530 650 540 654
rect 526 647 527 650
rect 529 647 540 650
rect 462 637 463 640
rect 465 637 473 640
rect 475 637 477 640
rect 489 639 495 645
rect 485 633 495 639
rect 530 645 540 647
rect 543 658 585 675
rect 543 657 563 658
rect 543 645 553 657
rect 558 656 561 657
rect 558 653 561 654
rect 569 654 585 658
rect 575 650 585 654
rect 571 647 572 650
rect 574 647 585 650
rect 507 637 508 640
rect 510 637 518 640
rect 520 637 522 640
rect 534 639 540 645
rect 530 633 540 639
rect 575 645 585 647
rect 588 658 630 675
rect 588 657 608 658
rect 588 645 598 657
rect 603 656 606 657
rect 603 653 606 654
rect 614 654 630 658
rect 620 650 630 654
rect 616 647 617 650
rect 619 647 630 650
rect 552 637 553 640
rect 555 637 563 640
rect 565 637 567 640
rect 579 639 585 645
rect 575 633 585 639
rect 620 645 630 647
rect 633 658 675 675
rect 633 657 653 658
rect 633 645 643 657
rect 648 656 651 657
rect 648 653 651 654
rect 659 654 675 658
rect 665 650 675 654
rect 661 647 662 650
rect 664 647 675 650
rect 597 637 598 640
rect 600 637 608 640
rect 610 637 612 640
rect 624 639 630 645
rect 620 633 630 639
rect 665 645 675 647
rect 678 658 720 675
rect 678 657 698 658
rect 678 645 688 657
rect 693 656 696 657
rect 693 653 696 654
rect 704 654 720 658
rect 710 650 720 654
rect 706 647 707 650
rect 709 647 720 650
rect 642 637 643 640
rect 645 637 653 640
rect 655 637 657 640
rect 669 639 675 645
rect 665 633 675 639
rect 710 645 720 647
rect 723 658 765 675
rect 723 657 743 658
rect 723 645 733 657
rect 738 656 741 657
rect 738 653 741 654
rect 749 654 765 658
rect 755 650 765 654
rect 751 647 752 650
rect 754 647 765 650
rect 687 637 688 640
rect 690 637 698 640
rect 700 637 702 640
rect 714 639 720 645
rect 710 633 720 639
rect 755 645 765 647
rect 768 658 810 675
rect 768 657 788 658
rect 768 645 778 657
rect 783 656 786 657
rect 783 653 786 654
rect 794 654 810 658
rect 800 650 810 654
rect 796 647 797 650
rect 799 647 810 650
rect 732 637 733 640
rect 735 637 743 640
rect 745 637 747 640
rect 759 639 765 645
rect 755 633 765 639
rect 800 645 810 647
rect 813 658 855 675
rect 813 657 833 658
rect 813 645 823 657
rect 828 656 831 657
rect 828 653 831 654
rect 839 654 855 658
rect 845 650 855 654
rect 841 647 842 650
rect 844 647 855 650
rect 777 637 778 640
rect 780 637 788 640
rect 790 637 792 640
rect 804 639 810 645
rect 800 633 810 639
rect 845 645 855 647
rect 858 658 900 675
rect 858 657 878 658
rect 858 645 868 657
rect 873 656 876 657
rect 873 653 876 654
rect 884 654 900 658
rect 890 650 900 654
rect 886 647 887 650
rect 889 647 900 650
rect 822 637 823 640
rect 825 637 833 640
rect 835 637 837 640
rect 849 639 855 645
rect 845 633 855 639
rect 890 645 900 647
rect 867 637 868 640
rect 870 637 878 640
rect 880 637 882 640
rect 894 639 900 645
rect 890 633 900 639
rect 3 613 45 630
rect 3 612 23 613
rect 3 600 13 612
rect 18 611 21 612
rect 18 608 21 609
rect 29 609 45 613
rect 35 605 45 609
rect 31 602 32 605
rect 34 602 45 605
rect 35 600 45 602
rect 48 613 90 630
rect 48 612 68 613
rect 48 600 58 612
rect 63 611 66 612
rect 63 608 66 609
rect 74 609 90 613
rect 80 605 90 609
rect 76 602 77 605
rect 79 602 90 605
rect 12 592 13 595
rect 15 592 23 595
rect 25 592 27 595
rect 39 594 45 600
rect 35 588 45 594
rect 80 600 90 602
rect 93 613 135 630
rect 93 612 113 613
rect 93 600 103 612
rect 108 611 111 612
rect 108 608 111 609
rect 119 609 135 613
rect 125 605 135 609
rect 121 602 122 605
rect 124 602 135 605
rect 57 592 58 595
rect 60 592 68 595
rect 70 592 72 595
rect 84 594 90 600
rect 80 588 90 594
rect 125 600 135 602
rect 138 613 180 630
rect 138 612 158 613
rect 138 600 148 612
rect 153 611 156 612
rect 153 608 156 609
rect 164 609 180 613
rect 170 605 180 609
rect 166 602 167 605
rect 169 602 180 605
rect 102 592 103 595
rect 105 592 113 595
rect 115 592 117 595
rect 129 594 135 600
rect 125 588 135 594
rect 170 600 180 602
rect 183 613 225 630
rect 183 612 203 613
rect 183 600 193 612
rect 198 611 201 612
rect 198 608 201 609
rect 209 609 225 613
rect 215 605 225 609
rect 211 602 212 605
rect 214 602 225 605
rect 147 592 148 595
rect 150 592 158 595
rect 160 592 162 595
rect 174 594 180 600
rect 170 588 180 594
rect 215 600 225 602
rect 228 613 270 630
rect 228 612 248 613
rect 228 600 238 612
rect 243 611 246 612
rect 243 608 246 609
rect 254 609 270 613
rect 260 605 270 609
rect 256 602 257 605
rect 259 602 270 605
rect 192 592 193 595
rect 195 592 203 595
rect 205 592 207 595
rect 219 594 225 600
rect 215 588 225 594
rect 260 600 270 602
rect 273 613 315 630
rect 273 612 293 613
rect 273 600 283 612
rect 288 611 291 612
rect 288 608 291 609
rect 299 609 315 613
rect 305 605 315 609
rect 301 602 302 605
rect 304 602 315 605
rect 237 592 238 595
rect 240 592 248 595
rect 250 592 252 595
rect 264 594 270 600
rect 260 588 270 594
rect 305 600 315 602
rect 318 613 360 630
rect 318 612 338 613
rect 318 600 328 612
rect 333 611 336 612
rect 333 608 336 609
rect 344 609 360 613
rect 350 605 360 609
rect 346 602 347 605
rect 349 602 360 605
rect 282 592 283 595
rect 285 592 293 595
rect 295 592 297 595
rect 309 594 315 600
rect 305 588 315 594
rect 350 600 360 602
rect 363 613 405 630
rect 363 612 383 613
rect 363 600 373 612
rect 378 611 381 612
rect 378 608 381 609
rect 389 609 405 613
rect 395 605 405 609
rect 391 602 392 605
rect 394 602 405 605
rect 327 592 328 595
rect 330 592 338 595
rect 340 592 342 595
rect 354 594 360 600
rect 350 588 360 594
rect 395 600 405 602
rect 408 613 450 630
rect 408 612 428 613
rect 408 600 418 612
rect 423 611 426 612
rect 423 608 426 609
rect 434 609 450 613
rect 440 605 450 609
rect 436 602 437 605
rect 439 602 450 605
rect 372 592 373 595
rect 375 592 383 595
rect 385 592 387 595
rect 399 594 405 600
rect 395 588 405 594
rect 440 600 450 602
rect 453 613 495 630
rect 453 612 473 613
rect 453 600 463 612
rect 468 611 471 612
rect 468 608 471 609
rect 479 609 495 613
rect 485 605 495 609
rect 481 602 482 605
rect 484 602 495 605
rect 417 592 418 595
rect 420 592 428 595
rect 430 592 432 595
rect 444 594 450 600
rect 440 588 450 594
rect 485 600 495 602
rect 498 613 540 630
rect 498 612 518 613
rect 498 600 508 612
rect 513 611 516 612
rect 513 608 516 609
rect 524 609 540 613
rect 530 605 540 609
rect 526 602 527 605
rect 529 602 540 605
rect 462 592 463 595
rect 465 592 473 595
rect 475 592 477 595
rect 489 594 495 600
rect 485 588 495 594
rect 530 600 540 602
rect 543 613 585 630
rect 543 612 563 613
rect 543 600 553 612
rect 558 611 561 612
rect 558 608 561 609
rect 569 609 585 613
rect 575 605 585 609
rect 571 602 572 605
rect 574 602 585 605
rect 507 592 508 595
rect 510 592 518 595
rect 520 592 522 595
rect 534 594 540 600
rect 530 588 540 594
rect 575 600 585 602
rect 588 613 630 630
rect 588 612 608 613
rect 588 600 598 612
rect 603 611 606 612
rect 603 608 606 609
rect 614 609 630 613
rect 620 605 630 609
rect 616 602 617 605
rect 619 602 630 605
rect 552 592 553 595
rect 555 592 563 595
rect 565 592 567 595
rect 579 594 585 600
rect 575 588 585 594
rect 620 600 630 602
rect 633 613 675 630
rect 633 612 653 613
rect 633 600 643 612
rect 648 611 651 612
rect 648 608 651 609
rect 659 609 675 613
rect 665 605 675 609
rect 661 602 662 605
rect 664 602 675 605
rect 597 592 598 595
rect 600 592 608 595
rect 610 592 612 595
rect 624 594 630 600
rect 620 588 630 594
rect 665 600 675 602
rect 678 613 720 630
rect 678 612 698 613
rect 678 600 688 612
rect 693 611 696 612
rect 693 608 696 609
rect 704 609 720 613
rect 710 605 720 609
rect 706 602 707 605
rect 709 602 720 605
rect 642 592 643 595
rect 645 592 653 595
rect 655 592 657 595
rect 669 594 675 600
rect 665 588 675 594
rect 710 600 720 602
rect 723 613 765 630
rect 723 612 743 613
rect 723 600 733 612
rect 738 611 741 612
rect 738 608 741 609
rect 749 609 765 613
rect 755 605 765 609
rect 751 602 752 605
rect 754 602 765 605
rect 687 592 688 595
rect 690 592 698 595
rect 700 592 702 595
rect 714 594 720 600
rect 710 588 720 594
rect 755 600 765 602
rect 768 613 810 630
rect 768 612 788 613
rect 768 600 778 612
rect 783 611 786 612
rect 783 608 786 609
rect 794 609 810 613
rect 800 605 810 609
rect 796 602 797 605
rect 799 602 810 605
rect 732 592 733 595
rect 735 592 743 595
rect 745 592 747 595
rect 759 594 765 600
rect 755 588 765 594
rect 800 600 810 602
rect 813 613 855 630
rect 813 612 833 613
rect 813 600 823 612
rect 828 611 831 612
rect 828 608 831 609
rect 839 609 855 613
rect 845 605 855 609
rect 841 602 842 605
rect 844 602 855 605
rect 777 592 778 595
rect 780 592 788 595
rect 790 592 792 595
rect 804 594 810 600
rect 800 588 810 594
rect 845 600 855 602
rect 858 613 900 630
rect 858 612 878 613
rect 858 600 868 612
rect 873 611 876 612
rect 873 608 876 609
rect 884 609 900 613
rect 890 605 900 609
rect 886 602 887 605
rect 889 602 900 605
rect 822 592 823 595
rect 825 592 833 595
rect 835 592 837 595
rect 849 594 855 600
rect 845 588 855 594
rect 890 600 900 602
rect 867 592 868 595
rect 870 592 878 595
rect 880 592 882 595
rect 894 594 900 600
rect 890 588 900 594
rect 3 568 45 585
rect 3 567 23 568
rect 3 555 13 567
rect 18 566 21 567
rect 18 563 21 564
rect 29 564 45 568
rect 35 560 45 564
rect 31 557 32 560
rect 34 557 45 560
rect 35 555 45 557
rect 48 568 90 585
rect 48 567 68 568
rect 48 555 58 567
rect 63 566 66 567
rect 63 563 66 564
rect 74 564 90 568
rect 80 560 90 564
rect 76 557 77 560
rect 79 557 90 560
rect 12 547 13 550
rect 15 547 23 550
rect 25 547 27 550
rect 39 549 45 555
rect 35 543 45 549
rect 80 555 90 557
rect 93 568 135 585
rect 93 567 113 568
rect 93 555 103 567
rect 108 566 111 567
rect 108 563 111 564
rect 119 564 135 568
rect 125 560 135 564
rect 121 557 122 560
rect 124 557 135 560
rect 57 547 58 550
rect 60 547 68 550
rect 70 547 72 550
rect 84 549 90 555
rect 80 543 90 549
rect 125 555 135 557
rect 138 568 180 585
rect 138 567 158 568
rect 138 555 148 567
rect 153 566 156 567
rect 153 563 156 564
rect 164 564 180 568
rect 170 560 180 564
rect 166 557 167 560
rect 169 557 180 560
rect 102 547 103 550
rect 105 547 113 550
rect 115 547 117 550
rect 129 549 135 555
rect 125 543 135 549
rect 170 555 180 557
rect 183 568 225 585
rect 183 567 203 568
rect 183 555 193 567
rect 198 566 201 567
rect 198 563 201 564
rect 209 564 225 568
rect 215 560 225 564
rect 211 557 212 560
rect 214 557 225 560
rect 147 547 148 550
rect 150 547 158 550
rect 160 547 162 550
rect 174 549 180 555
rect 170 543 180 549
rect 215 555 225 557
rect 228 568 270 585
rect 228 567 248 568
rect 228 555 238 567
rect 243 566 246 567
rect 243 563 246 564
rect 254 564 270 568
rect 260 560 270 564
rect 256 557 257 560
rect 259 557 270 560
rect 192 547 193 550
rect 195 547 203 550
rect 205 547 207 550
rect 219 549 225 555
rect 215 543 225 549
rect 260 555 270 557
rect 273 568 315 585
rect 273 567 293 568
rect 273 555 283 567
rect 288 566 291 567
rect 288 563 291 564
rect 299 564 315 568
rect 305 560 315 564
rect 301 557 302 560
rect 304 557 315 560
rect 237 547 238 550
rect 240 547 248 550
rect 250 547 252 550
rect 264 549 270 555
rect 260 543 270 549
rect 305 555 315 557
rect 318 568 360 585
rect 318 567 338 568
rect 318 555 328 567
rect 333 566 336 567
rect 333 563 336 564
rect 344 564 360 568
rect 350 560 360 564
rect 346 557 347 560
rect 349 557 360 560
rect 282 547 283 550
rect 285 547 293 550
rect 295 547 297 550
rect 309 549 315 555
rect 305 543 315 549
rect 350 555 360 557
rect 363 568 405 585
rect 363 567 383 568
rect 363 555 373 567
rect 378 566 381 567
rect 378 563 381 564
rect 389 564 405 568
rect 395 560 405 564
rect 391 557 392 560
rect 394 557 405 560
rect 327 547 328 550
rect 330 547 338 550
rect 340 547 342 550
rect 354 549 360 555
rect 350 543 360 549
rect 395 555 405 557
rect 408 568 450 585
rect 408 567 428 568
rect 408 555 418 567
rect 423 566 426 567
rect 423 563 426 564
rect 434 564 450 568
rect 440 560 450 564
rect 436 557 437 560
rect 439 557 450 560
rect 372 547 373 550
rect 375 547 383 550
rect 385 547 387 550
rect 399 549 405 555
rect 395 543 405 549
rect 440 555 450 557
rect 453 568 495 585
rect 453 567 473 568
rect 453 555 463 567
rect 468 566 471 567
rect 468 563 471 564
rect 479 564 495 568
rect 485 560 495 564
rect 481 557 482 560
rect 484 557 495 560
rect 417 547 418 550
rect 420 547 428 550
rect 430 547 432 550
rect 444 549 450 555
rect 440 543 450 549
rect 485 555 495 557
rect 498 568 540 585
rect 498 567 518 568
rect 498 555 508 567
rect 513 566 516 567
rect 513 563 516 564
rect 524 564 540 568
rect 530 560 540 564
rect 526 557 527 560
rect 529 557 540 560
rect 462 547 463 550
rect 465 547 473 550
rect 475 547 477 550
rect 489 549 495 555
rect 485 543 495 549
rect 530 555 540 557
rect 543 568 585 585
rect 543 567 563 568
rect 543 555 553 567
rect 558 566 561 567
rect 558 563 561 564
rect 569 564 585 568
rect 575 560 585 564
rect 571 557 572 560
rect 574 557 585 560
rect 507 547 508 550
rect 510 547 518 550
rect 520 547 522 550
rect 534 549 540 555
rect 530 543 540 549
rect 575 555 585 557
rect 588 568 630 585
rect 588 567 608 568
rect 588 555 598 567
rect 603 566 606 567
rect 603 563 606 564
rect 614 564 630 568
rect 620 560 630 564
rect 616 557 617 560
rect 619 557 630 560
rect 552 547 553 550
rect 555 547 563 550
rect 565 547 567 550
rect 579 549 585 555
rect 575 543 585 549
rect 620 555 630 557
rect 633 568 675 585
rect 633 567 653 568
rect 633 555 643 567
rect 648 566 651 567
rect 648 563 651 564
rect 659 564 675 568
rect 665 560 675 564
rect 661 557 662 560
rect 664 557 675 560
rect 597 547 598 550
rect 600 547 608 550
rect 610 547 612 550
rect 624 549 630 555
rect 620 543 630 549
rect 665 555 675 557
rect 678 568 720 585
rect 678 567 698 568
rect 678 555 688 567
rect 693 566 696 567
rect 693 563 696 564
rect 704 564 720 568
rect 710 560 720 564
rect 706 557 707 560
rect 709 557 720 560
rect 642 547 643 550
rect 645 547 653 550
rect 655 547 657 550
rect 669 549 675 555
rect 665 543 675 549
rect 710 555 720 557
rect 723 568 765 585
rect 723 567 743 568
rect 723 555 733 567
rect 738 566 741 567
rect 738 563 741 564
rect 749 564 765 568
rect 755 560 765 564
rect 751 557 752 560
rect 754 557 765 560
rect 687 547 688 550
rect 690 547 698 550
rect 700 547 702 550
rect 714 549 720 555
rect 710 543 720 549
rect 755 555 765 557
rect 768 568 810 585
rect 768 567 788 568
rect 768 555 778 567
rect 783 566 786 567
rect 783 563 786 564
rect 794 564 810 568
rect 800 560 810 564
rect 796 557 797 560
rect 799 557 810 560
rect 732 547 733 550
rect 735 547 743 550
rect 745 547 747 550
rect 759 549 765 555
rect 755 543 765 549
rect 800 555 810 557
rect 813 568 855 585
rect 813 567 833 568
rect 813 555 823 567
rect 828 566 831 567
rect 828 563 831 564
rect 839 564 855 568
rect 845 560 855 564
rect 841 557 842 560
rect 844 557 855 560
rect 777 547 778 550
rect 780 547 788 550
rect 790 547 792 550
rect 804 549 810 555
rect 800 543 810 549
rect 845 555 855 557
rect 858 568 900 585
rect 858 567 878 568
rect 858 555 868 567
rect 873 566 876 567
rect 873 563 876 564
rect 884 564 900 568
rect 890 560 900 564
rect 886 557 887 560
rect 889 557 900 560
rect 822 547 823 550
rect 825 547 833 550
rect 835 547 837 550
rect 849 549 855 555
rect 845 543 855 549
rect 890 555 900 557
rect 867 547 868 550
rect 870 547 878 550
rect 880 547 882 550
rect 894 549 900 555
rect 890 543 900 549
rect 3 523 45 540
rect 3 522 23 523
rect 3 510 13 522
rect 18 521 21 522
rect 18 518 21 519
rect 29 519 45 523
rect 35 515 45 519
rect 31 512 32 515
rect 34 512 45 515
rect 35 510 45 512
rect 48 523 90 540
rect 48 522 68 523
rect 48 510 58 522
rect 63 521 66 522
rect 63 518 66 519
rect 74 519 90 523
rect 80 515 90 519
rect 76 512 77 515
rect 79 512 90 515
rect 12 502 13 505
rect 15 502 23 505
rect 25 502 27 505
rect 39 504 45 510
rect 35 498 45 504
rect 80 510 90 512
rect 93 523 135 540
rect 93 522 113 523
rect 93 510 103 522
rect 108 521 111 522
rect 108 518 111 519
rect 119 519 135 523
rect 125 515 135 519
rect 121 512 122 515
rect 124 512 135 515
rect 57 502 58 505
rect 60 502 68 505
rect 70 502 72 505
rect 84 504 90 510
rect 80 498 90 504
rect 125 510 135 512
rect 138 523 180 540
rect 138 522 158 523
rect 138 510 148 522
rect 153 521 156 522
rect 153 518 156 519
rect 164 519 180 523
rect 170 515 180 519
rect 166 512 167 515
rect 169 512 180 515
rect 102 502 103 505
rect 105 502 113 505
rect 115 502 117 505
rect 129 504 135 510
rect 125 498 135 504
rect 170 510 180 512
rect 183 523 225 540
rect 183 522 203 523
rect 183 510 193 522
rect 198 521 201 522
rect 198 518 201 519
rect 209 519 225 523
rect 215 515 225 519
rect 211 512 212 515
rect 214 512 225 515
rect 147 502 148 505
rect 150 502 158 505
rect 160 502 162 505
rect 174 504 180 510
rect 170 498 180 504
rect 215 510 225 512
rect 228 523 270 540
rect 228 522 248 523
rect 228 510 238 522
rect 243 521 246 522
rect 243 518 246 519
rect 254 519 270 523
rect 260 515 270 519
rect 256 512 257 515
rect 259 512 270 515
rect 192 502 193 505
rect 195 502 203 505
rect 205 502 207 505
rect 219 504 225 510
rect 215 498 225 504
rect 260 510 270 512
rect 273 523 315 540
rect 273 522 293 523
rect 273 510 283 522
rect 288 521 291 522
rect 288 518 291 519
rect 299 519 315 523
rect 305 515 315 519
rect 301 512 302 515
rect 304 512 315 515
rect 237 502 238 505
rect 240 502 248 505
rect 250 502 252 505
rect 264 504 270 510
rect 260 498 270 504
rect 305 510 315 512
rect 318 523 360 540
rect 318 522 338 523
rect 318 510 328 522
rect 333 521 336 522
rect 333 518 336 519
rect 344 519 360 523
rect 350 515 360 519
rect 346 512 347 515
rect 349 512 360 515
rect 282 502 283 505
rect 285 502 293 505
rect 295 502 297 505
rect 309 504 315 510
rect 305 498 315 504
rect 350 510 360 512
rect 363 523 405 540
rect 363 522 383 523
rect 363 510 373 522
rect 378 521 381 522
rect 378 518 381 519
rect 389 519 405 523
rect 395 515 405 519
rect 391 512 392 515
rect 394 512 405 515
rect 327 502 328 505
rect 330 502 338 505
rect 340 502 342 505
rect 354 504 360 510
rect 350 498 360 504
rect 395 510 405 512
rect 408 523 450 540
rect 408 522 428 523
rect 408 510 418 522
rect 423 521 426 522
rect 423 518 426 519
rect 434 519 450 523
rect 440 515 450 519
rect 436 512 437 515
rect 439 512 450 515
rect 372 502 373 505
rect 375 502 383 505
rect 385 502 387 505
rect 399 504 405 510
rect 395 498 405 504
rect 440 510 450 512
rect 453 523 495 540
rect 453 522 473 523
rect 453 510 463 522
rect 468 521 471 522
rect 468 518 471 519
rect 479 519 495 523
rect 485 515 495 519
rect 481 512 482 515
rect 484 512 495 515
rect 417 502 418 505
rect 420 502 428 505
rect 430 502 432 505
rect 444 504 450 510
rect 440 498 450 504
rect 485 510 495 512
rect 498 523 540 540
rect 498 522 518 523
rect 498 510 508 522
rect 513 521 516 522
rect 513 518 516 519
rect 524 519 540 523
rect 530 515 540 519
rect 526 512 527 515
rect 529 512 540 515
rect 462 502 463 505
rect 465 502 473 505
rect 475 502 477 505
rect 489 504 495 510
rect 485 498 495 504
rect 530 510 540 512
rect 543 523 585 540
rect 543 522 563 523
rect 543 510 553 522
rect 558 521 561 522
rect 558 518 561 519
rect 569 519 585 523
rect 575 515 585 519
rect 571 512 572 515
rect 574 512 585 515
rect 507 502 508 505
rect 510 502 518 505
rect 520 502 522 505
rect 534 504 540 510
rect 530 498 540 504
rect 575 510 585 512
rect 588 523 630 540
rect 588 522 608 523
rect 588 510 598 522
rect 603 521 606 522
rect 603 518 606 519
rect 614 519 630 523
rect 620 515 630 519
rect 616 512 617 515
rect 619 512 630 515
rect 552 502 553 505
rect 555 502 563 505
rect 565 502 567 505
rect 579 504 585 510
rect 575 498 585 504
rect 620 510 630 512
rect 633 523 675 540
rect 633 522 653 523
rect 633 510 643 522
rect 648 521 651 522
rect 648 518 651 519
rect 659 519 675 523
rect 665 515 675 519
rect 661 512 662 515
rect 664 512 675 515
rect 597 502 598 505
rect 600 502 608 505
rect 610 502 612 505
rect 624 504 630 510
rect 620 498 630 504
rect 665 510 675 512
rect 678 523 720 540
rect 678 522 698 523
rect 678 510 688 522
rect 693 521 696 522
rect 693 518 696 519
rect 704 519 720 523
rect 710 515 720 519
rect 706 512 707 515
rect 709 512 720 515
rect 642 502 643 505
rect 645 502 653 505
rect 655 502 657 505
rect 669 504 675 510
rect 665 498 675 504
rect 710 510 720 512
rect 723 523 765 540
rect 723 522 743 523
rect 723 510 733 522
rect 738 521 741 522
rect 738 518 741 519
rect 749 519 765 523
rect 755 515 765 519
rect 751 512 752 515
rect 754 512 765 515
rect 687 502 688 505
rect 690 502 698 505
rect 700 502 702 505
rect 714 504 720 510
rect 710 498 720 504
rect 755 510 765 512
rect 768 523 810 540
rect 768 522 788 523
rect 768 510 778 522
rect 783 521 786 522
rect 783 518 786 519
rect 794 519 810 523
rect 800 515 810 519
rect 796 512 797 515
rect 799 512 810 515
rect 732 502 733 505
rect 735 502 743 505
rect 745 502 747 505
rect 759 504 765 510
rect 755 498 765 504
rect 800 510 810 512
rect 813 523 855 540
rect 813 522 833 523
rect 813 510 823 522
rect 828 521 831 522
rect 828 518 831 519
rect 839 519 855 523
rect 845 515 855 519
rect 841 512 842 515
rect 844 512 855 515
rect 777 502 778 505
rect 780 502 788 505
rect 790 502 792 505
rect 804 504 810 510
rect 800 498 810 504
rect 845 510 855 512
rect 858 523 900 540
rect 858 522 878 523
rect 858 510 868 522
rect 873 521 876 522
rect 873 518 876 519
rect 884 519 900 523
rect 890 515 900 519
rect 886 512 887 515
rect 889 512 900 515
rect 822 502 823 505
rect 825 502 833 505
rect 835 502 837 505
rect 849 504 855 510
rect 845 498 855 504
rect 890 510 900 512
rect 867 502 868 505
rect 870 502 878 505
rect 880 502 882 505
rect 894 504 900 510
rect 890 498 900 504
rect 3 478 45 495
rect 3 477 23 478
rect 3 465 13 477
rect 18 476 21 477
rect 18 473 21 474
rect 29 474 45 478
rect 35 470 45 474
rect 31 467 32 470
rect 34 467 45 470
rect 35 465 45 467
rect 48 478 90 495
rect 48 477 68 478
rect 48 465 58 477
rect 63 476 66 477
rect 63 473 66 474
rect 74 474 90 478
rect 80 470 90 474
rect 76 467 77 470
rect 79 467 90 470
rect 12 457 13 460
rect 15 457 23 460
rect 25 457 27 460
rect 39 459 45 465
rect 35 453 45 459
rect 80 465 90 467
rect 93 478 135 495
rect 93 477 113 478
rect 93 465 103 477
rect 108 476 111 477
rect 108 473 111 474
rect 119 474 135 478
rect 125 470 135 474
rect 121 467 122 470
rect 124 467 135 470
rect 57 457 58 460
rect 60 457 68 460
rect 70 457 72 460
rect 84 459 90 465
rect 80 453 90 459
rect 125 465 135 467
rect 138 478 180 495
rect 138 477 158 478
rect 138 465 148 477
rect 153 476 156 477
rect 153 473 156 474
rect 164 474 180 478
rect 170 470 180 474
rect 166 467 167 470
rect 169 467 180 470
rect 102 457 103 460
rect 105 457 113 460
rect 115 457 117 460
rect 129 459 135 465
rect 125 453 135 459
rect 170 465 180 467
rect 183 478 225 495
rect 183 477 203 478
rect 183 465 193 477
rect 198 476 201 477
rect 198 473 201 474
rect 209 474 225 478
rect 215 470 225 474
rect 211 467 212 470
rect 214 467 225 470
rect 147 457 148 460
rect 150 457 158 460
rect 160 457 162 460
rect 174 459 180 465
rect 170 453 180 459
rect 215 465 225 467
rect 228 478 270 495
rect 228 477 248 478
rect 228 465 238 477
rect 243 476 246 477
rect 243 473 246 474
rect 254 474 270 478
rect 260 470 270 474
rect 256 467 257 470
rect 259 467 270 470
rect 192 457 193 460
rect 195 457 203 460
rect 205 457 207 460
rect 219 459 225 465
rect 215 453 225 459
rect 260 465 270 467
rect 273 478 315 495
rect 273 477 293 478
rect 273 465 283 477
rect 288 476 291 477
rect 288 473 291 474
rect 299 474 315 478
rect 305 470 315 474
rect 301 467 302 470
rect 304 467 315 470
rect 237 457 238 460
rect 240 457 248 460
rect 250 457 252 460
rect 264 459 270 465
rect 260 453 270 459
rect 305 465 315 467
rect 318 478 360 495
rect 318 477 338 478
rect 318 465 328 477
rect 333 476 336 477
rect 333 473 336 474
rect 344 474 360 478
rect 350 470 360 474
rect 346 467 347 470
rect 349 467 360 470
rect 282 457 283 460
rect 285 457 293 460
rect 295 457 297 460
rect 309 459 315 465
rect 305 453 315 459
rect 350 465 360 467
rect 363 478 405 495
rect 363 477 383 478
rect 363 465 373 477
rect 378 476 381 477
rect 378 473 381 474
rect 389 474 405 478
rect 395 470 405 474
rect 391 467 392 470
rect 394 467 405 470
rect 327 457 328 460
rect 330 457 338 460
rect 340 457 342 460
rect 354 459 360 465
rect 350 453 360 459
rect 395 465 405 467
rect 408 478 450 495
rect 408 477 428 478
rect 408 465 418 477
rect 423 476 426 477
rect 423 473 426 474
rect 434 474 450 478
rect 440 470 450 474
rect 436 467 437 470
rect 439 467 450 470
rect 372 457 373 460
rect 375 457 383 460
rect 385 457 387 460
rect 399 459 405 465
rect 395 453 405 459
rect 440 465 450 467
rect 453 478 495 495
rect 453 477 473 478
rect 453 465 463 477
rect 468 476 471 477
rect 468 473 471 474
rect 479 474 495 478
rect 485 470 495 474
rect 481 467 482 470
rect 484 467 495 470
rect 417 457 418 460
rect 420 457 428 460
rect 430 457 432 460
rect 444 459 450 465
rect 440 453 450 459
rect 485 465 495 467
rect 498 478 540 495
rect 498 477 518 478
rect 498 465 508 477
rect 513 476 516 477
rect 513 473 516 474
rect 524 474 540 478
rect 530 470 540 474
rect 526 467 527 470
rect 529 467 540 470
rect 462 457 463 460
rect 465 457 473 460
rect 475 457 477 460
rect 489 459 495 465
rect 485 453 495 459
rect 530 465 540 467
rect 543 478 585 495
rect 543 477 563 478
rect 543 465 553 477
rect 558 476 561 477
rect 558 473 561 474
rect 569 474 585 478
rect 575 470 585 474
rect 571 467 572 470
rect 574 467 585 470
rect 507 457 508 460
rect 510 457 518 460
rect 520 457 522 460
rect 534 459 540 465
rect 530 453 540 459
rect 575 465 585 467
rect 588 478 630 495
rect 588 477 608 478
rect 588 465 598 477
rect 603 476 606 477
rect 603 473 606 474
rect 614 474 630 478
rect 620 470 630 474
rect 616 467 617 470
rect 619 467 630 470
rect 552 457 553 460
rect 555 457 563 460
rect 565 457 567 460
rect 579 459 585 465
rect 575 453 585 459
rect 620 465 630 467
rect 633 478 675 495
rect 633 477 653 478
rect 633 465 643 477
rect 648 476 651 477
rect 648 473 651 474
rect 659 474 675 478
rect 665 470 675 474
rect 661 467 662 470
rect 664 467 675 470
rect 597 457 598 460
rect 600 457 608 460
rect 610 457 612 460
rect 624 459 630 465
rect 620 453 630 459
rect 665 465 675 467
rect 678 478 720 495
rect 678 477 698 478
rect 678 465 688 477
rect 693 476 696 477
rect 693 473 696 474
rect 704 474 720 478
rect 710 470 720 474
rect 706 467 707 470
rect 709 467 720 470
rect 642 457 643 460
rect 645 457 653 460
rect 655 457 657 460
rect 669 459 675 465
rect 665 453 675 459
rect 710 465 720 467
rect 723 478 765 495
rect 723 477 743 478
rect 723 465 733 477
rect 738 476 741 477
rect 738 473 741 474
rect 749 474 765 478
rect 755 470 765 474
rect 751 467 752 470
rect 754 467 765 470
rect 687 457 688 460
rect 690 457 698 460
rect 700 457 702 460
rect 714 459 720 465
rect 710 453 720 459
rect 755 465 765 467
rect 768 478 810 495
rect 768 477 788 478
rect 768 465 778 477
rect 783 476 786 477
rect 783 473 786 474
rect 794 474 810 478
rect 800 470 810 474
rect 796 467 797 470
rect 799 467 810 470
rect 732 457 733 460
rect 735 457 743 460
rect 745 457 747 460
rect 759 459 765 465
rect 755 453 765 459
rect 800 465 810 467
rect 813 478 855 495
rect 813 477 833 478
rect 813 465 823 477
rect 828 476 831 477
rect 828 473 831 474
rect 839 474 855 478
rect 845 470 855 474
rect 841 467 842 470
rect 844 467 855 470
rect 777 457 778 460
rect 780 457 788 460
rect 790 457 792 460
rect 804 459 810 465
rect 800 453 810 459
rect 845 465 855 467
rect 858 478 900 495
rect 858 477 878 478
rect 858 465 868 477
rect 873 476 876 477
rect 873 473 876 474
rect 884 474 900 478
rect 890 470 900 474
rect 886 467 887 470
rect 889 467 900 470
rect 822 457 823 460
rect 825 457 833 460
rect 835 457 837 460
rect 849 459 855 465
rect 845 453 855 459
rect 890 465 900 467
rect 867 457 868 460
rect 870 457 878 460
rect 880 457 882 460
rect 894 459 900 465
rect 890 453 900 459
rect 3 433 45 450
rect 3 432 23 433
rect 3 420 13 432
rect 18 431 21 432
rect 18 428 21 429
rect 29 429 45 433
rect 35 425 45 429
rect 31 422 32 425
rect 34 422 45 425
rect 35 420 45 422
rect 48 433 90 450
rect 48 432 68 433
rect 48 420 58 432
rect 63 431 66 432
rect 63 428 66 429
rect 74 429 90 433
rect 80 425 90 429
rect 76 422 77 425
rect 79 422 90 425
rect 12 412 13 415
rect 15 412 23 415
rect 25 412 27 415
rect 39 414 45 420
rect 35 408 45 414
rect 80 420 90 422
rect 93 433 135 450
rect 93 432 113 433
rect 93 420 103 432
rect 108 431 111 432
rect 108 428 111 429
rect 119 429 135 433
rect 125 425 135 429
rect 121 422 122 425
rect 124 422 135 425
rect 57 412 58 415
rect 60 412 68 415
rect 70 412 72 415
rect 84 414 90 420
rect 80 408 90 414
rect 125 420 135 422
rect 138 433 180 450
rect 138 432 158 433
rect 138 420 148 432
rect 153 431 156 432
rect 153 428 156 429
rect 164 429 180 433
rect 170 425 180 429
rect 166 422 167 425
rect 169 422 180 425
rect 102 412 103 415
rect 105 412 113 415
rect 115 412 117 415
rect 129 414 135 420
rect 125 408 135 414
rect 170 420 180 422
rect 183 433 225 450
rect 183 432 203 433
rect 183 420 193 432
rect 198 431 201 432
rect 198 428 201 429
rect 209 429 225 433
rect 215 425 225 429
rect 211 422 212 425
rect 214 422 225 425
rect 147 412 148 415
rect 150 412 158 415
rect 160 412 162 415
rect 174 414 180 420
rect 170 408 180 414
rect 215 420 225 422
rect 228 433 270 450
rect 228 432 248 433
rect 228 420 238 432
rect 243 431 246 432
rect 243 428 246 429
rect 254 429 270 433
rect 260 425 270 429
rect 256 422 257 425
rect 259 422 270 425
rect 192 412 193 415
rect 195 412 203 415
rect 205 412 207 415
rect 219 414 225 420
rect 215 408 225 414
rect 260 420 270 422
rect 273 433 315 450
rect 273 432 293 433
rect 273 420 283 432
rect 288 431 291 432
rect 288 428 291 429
rect 299 429 315 433
rect 305 425 315 429
rect 301 422 302 425
rect 304 422 315 425
rect 237 412 238 415
rect 240 412 248 415
rect 250 412 252 415
rect 264 414 270 420
rect 260 408 270 414
rect 305 420 315 422
rect 318 433 360 450
rect 318 432 338 433
rect 318 420 328 432
rect 333 431 336 432
rect 333 428 336 429
rect 344 429 360 433
rect 350 425 360 429
rect 346 422 347 425
rect 349 422 360 425
rect 282 412 283 415
rect 285 412 293 415
rect 295 412 297 415
rect 309 414 315 420
rect 305 408 315 414
rect 350 420 360 422
rect 363 433 405 450
rect 363 432 383 433
rect 363 420 373 432
rect 378 431 381 432
rect 378 428 381 429
rect 389 429 405 433
rect 395 425 405 429
rect 391 422 392 425
rect 394 422 405 425
rect 327 412 328 415
rect 330 412 338 415
rect 340 412 342 415
rect 354 414 360 420
rect 350 408 360 414
rect 395 420 405 422
rect 408 433 450 450
rect 408 432 428 433
rect 408 420 418 432
rect 423 431 426 432
rect 423 428 426 429
rect 434 429 450 433
rect 440 425 450 429
rect 436 422 437 425
rect 439 422 450 425
rect 372 412 373 415
rect 375 412 383 415
rect 385 412 387 415
rect 399 414 405 420
rect 395 408 405 414
rect 440 420 450 422
rect 453 433 495 450
rect 453 432 473 433
rect 453 420 463 432
rect 468 431 471 432
rect 468 428 471 429
rect 479 429 495 433
rect 485 425 495 429
rect 481 422 482 425
rect 484 422 495 425
rect 417 412 418 415
rect 420 412 428 415
rect 430 412 432 415
rect 444 414 450 420
rect 440 408 450 414
rect 485 420 495 422
rect 498 433 540 450
rect 498 432 518 433
rect 498 420 508 432
rect 513 431 516 432
rect 513 428 516 429
rect 524 429 540 433
rect 530 425 540 429
rect 526 422 527 425
rect 529 422 540 425
rect 462 412 463 415
rect 465 412 473 415
rect 475 412 477 415
rect 489 414 495 420
rect 485 408 495 414
rect 530 420 540 422
rect 543 433 585 450
rect 543 432 563 433
rect 543 420 553 432
rect 558 431 561 432
rect 558 428 561 429
rect 569 429 585 433
rect 575 425 585 429
rect 571 422 572 425
rect 574 422 585 425
rect 507 412 508 415
rect 510 412 518 415
rect 520 412 522 415
rect 534 414 540 420
rect 530 408 540 414
rect 575 420 585 422
rect 588 433 630 450
rect 588 432 608 433
rect 588 420 598 432
rect 603 431 606 432
rect 603 428 606 429
rect 614 429 630 433
rect 620 425 630 429
rect 616 422 617 425
rect 619 422 630 425
rect 552 412 553 415
rect 555 412 563 415
rect 565 412 567 415
rect 579 414 585 420
rect 575 408 585 414
rect 620 420 630 422
rect 633 433 675 450
rect 633 432 653 433
rect 633 420 643 432
rect 648 431 651 432
rect 648 428 651 429
rect 659 429 675 433
rect 665 425 675 429
rect 661 422 662 425
rect 664 422 675 425
rect 597 412 598 415
rect 600 412 608 415
rect 610 412 612 415
rect 624 414 630 420
rect 620 408 630 414
rect 665 420 675 422
rect 678 433 720 450
rect 678 432 698 433
rect 678 420 688 432
rect 693 431 696 432
rect 693 428 696 429
rect 704 429 720 433
rect 710 425 720 429
rect 706 422 707 425
rect 709 422 720 425
rect 642 412 643 415
rect 645 412 653 415
rect 655 412 657 415
rect 669 414 675 420
rect 665 408 675 414
rect 710 420 720 422
rect 723 433 765 450
rect 723 432 743 433
rect 723 420 733 432
rect 738 431 741 432
rect 738 428 741 429
rect 749 429 765 433
rect 755 425 765 429
rect 751 422 752 425
rect 754 422 765 425
rect 687 412 688 415
rect 690 412 698 415
rect 700 412 702 415
rect 714 414 720 420
rect 710 408 720 414
rect 755 420 765 422
rect 768 433 810 450
rect 768 432 788 433
rect 768 420 778 432
rect 783 431 786 432
rect 783 428 786 429
rect 794 429 810 433
rect 800 425 810 429
rect 796 422 797 425
rect 799 422 810 425
rect 732 412 733 415
rect 735 412 743 415
rect 745 412 747 415
rect 759 414 765 420
rect 755 408 765 414
rect 800 420 810 422
rect 813 433 855 450
rect 813 432 833 433
rect 813 420 823 432
rect 828 431 831 432
rect 828 428 831 429
rect 839 429 855 433
rect 845 425 855 429
rect 841 422 842 425
rect 844 422 855 425
rect 777 412 778 415
rect 780 412 788 415
rect 790 412 792 415
rect 804 414 810 420
rect 800 408 810 414
rect 845 420 855 422
rect 858 433 900 450
rect 858 432 878 433
rect 858 420 868 432
rect 873 431 876 432
rect 873 428 876 429
rect 884 429 900 433
rect 890 425 900 429
rect 886 422 887 425
rect 889 422 900 425
rect 822 412 823 415
rect 825 412 833 415
rect 835 412 837 415
rect 849 414 855 420
rect 845 408 855 414
rect 890 420 900 422
rect 867 412 868 415
rect 870 412 878 415
rect 880 412 882 415
rect 894 414 900 420
rect 890 408 900 414
rect 3 388 45 405
rect 3 387 23 388
rect 3 375 13 387
rect 18 386 21 387
rect 18 383 21 384
rect 29 384 45 388
rect 35 380 45 384
rect 31 377 32 380
rect 34 377 45 380
rect 35 375 45 377
rect 48 388 90 405
rect 48 387 68 388
rect 48 375 58 387
rect 63 386 66 387
rect 63 383 66 384
rect 74 384 90 388
rect 80 380 90 384
rect 76 377 77 380
rect 79 377 90 380
rect 12 367 13 370
rect 15 367 23 370
rect 25 367 27 370
rect 39 369 45 375
rect 35 363 45 369
rect 80 375 90 377
rect 93 388 135 405
rect 93 387 113 388
rect 93 375 103 387
rect 108 386 111 387
rect 108 383 111 384
rect 119 384 135 388
rect 125 380 135 384
rect 121 377 122 380
rect 124 377 135 380
rect 57 367 58 370
rect 60 367 68 370
rect 70 367 72 370
rect 84 369 90 375
rect 80 363 90 369
rect 125 375 135 377
rect 138 388 180 405
rect 138 387 158 388
rect 138 375 148 387
rect 153 386 156 387
rect 153 383 156 384
rect 164 384 180 388
rect 170 380 180 384
rect 166 377 167 380
rect 169 377 180 380
rect 102 367 103 370
rect 105 367 113 370
rect 115 367 117 370
rect 129 369 135 375
rect 125 363 135 369
rect 170 375 180 377
rect 183 388 225 405
rect 183 387 203 388
rect 183 375 193 387
rect 198 386 201 387
rect 198 383 201 384
rect 209 384 225 388
rect 215 380 225 384
rect 211 377 212 380
rect 214 377 225 380
rect 147 367 148 370
rect 150 367 158 370
rect 160 367 162 370
rect 174 369 180 375
rect 170 363 180 369
rect 215 375 225 377
rect 228 388 270 405
rect 228 387 248 388
rect 228 375 238 387
rect 243 386 246 387
rect 243 383 246 384
rect 254 384 270 388
rect 260 380 270 384
rect 256 377 257 380
rect 259 377 270 380
rect 192 367 193 370
rect 195 367 203 370
rect 205 367 207 370
rect 219 369 225 375
rect 215 363 225 369
rect 260 375 270 377
rect 273 388 315 405
rect 273 387 293 388
rect 273 375 283 387
rect 288 386 291 387
rect 288 383 291 384
rect 299 384 315 388
rect 305 380 315 384
rect 301 377 302 380
rect 304 377 315 380
rect 237 367 238 370
rect 240 367 248 370
rect 250 367 252 370
rect 264 369 270 375
rect 260 363 270 369
rect 305 375 315 377
rect 318 388 360 405
rect 318 387 338 388
rect 318 375 328 387
rect 333 386 336 387
rect 333 383 336 384
rect 344 384 360 388
rect 350 380 360 384
rect 346 377 347 380
rect 349 377 360 380
rect 282 367 283 370
rect 285 367 293 370
rect 295 367 297 370
rect 309 369 315 375
rect 305 363 315 369
rect 350 375 360 377
rect 363 388 405 405
rect 363 387 383 388
rect 363 375 373 387
rect 378 386 381 387
rect 378 383 381 384
rect 389 384 405 388
rect 395 380 405 384
rect 391 377 392 380
rect 394 377 405 380
rect 327 367 328 370
rect 330 367 338 370
rect 340 367 342 370
rect 354 369 360 375
rect 350 363 360 369
rect 395 375 405 377
rect 408 388 450 405
rect 408 387 428 388
rect 408 375 418 387
rect 423 386 426 387
rect 423 383 426 384
rect 434 384 450 388
rect 440 380 450 384
rect 436 377 437 380
rect 439 377 450 380
rect 372 367 373 370
rect 375 367 383 370
rect 385 367 387 370
rect 399 369 405 375
rect 395 363 405 369
rect 440 375 450 377
rect 453 388 495 405
rect 453 387 473 388
rect 453 375 463 387
rect 468 386 471 387
rect 468 383 471 384
rect 479 384 495 388
rect 485 380 495 384
rect 481 377 482 380
rect 484 377 495 380
rect 417 367 418 370
rect 420 367 428 370
rect 430 367 432 370
rect 444 369 450 375
rect 440 363 450 369
rect 485 375 495 377
rect 498 388 540 405
rect 498 387 518 388
rect 498 375 508 387
rect 513 386 516 387
rect 513 383 516 384
rect 524 384 540 388
rect 530 380 540 384
rect 526 377 527 380
rect 529 377 540 380
rect 462 367 463 370
rect 465 367 473 370
rect 475 367 477 370
rect 489 369 495 375
rect 485 363 495 369
rect 530 375 540 377
rect 543 388 585 405
rect 543 387 563 388
rect 543 375 553 387
rect 558 386 561 387
rect 558 383 561 384
rect 569 384 585 388
rect 575 380 585 384
rect 571 377 572 380
rect 574 377 585 380
rect 507 367 508 370
rect 510 367 518 370
rect 520 367 522 370
rect 534 369 540 375
rect 530 363 540 369
rect 575 375 585 377
rect 588 388 630 405
rect 588 387 608 388
rect 588 375 598 387
rect 603 386 606 387
rect 603 383 606 384
rect 614 384 630 388
rect 620 380 630 384
rect 616 377 617 380
rect 619 377 630 380
rect 552 367 553 370
rect 555 367 563 370
rect 565 367 567 370
rect 579 369 585 375
rect 575 363 585 369
rect 620 375 630 377
rect 633 388 675 405
rect 633 387 653 388
rect 633 375 643 387
rect 648 386 651 387
rect 648 383 651 384
rect 659 384 675 388
rect 665 380 675 384
rect 661 377 662 380
rect 664 377 675 380
rect 597 367 598 370
rect 600 367 608 370
rect 610 367 612 370
rect 624 369 630 375
rect 620 363 630 369
rect 665 375 675 377
rect 678 388 720 405
rect 678 387 698 388
rect 678 375 688 387
rect 693 386 696 387
rect 693 383 696 384
rect 704 384 720 388
rect 710 380 720 384
rect 706 377 707 380
rect 709 377 720 380
rect 642 367 643 370
rect 645 367 653 370
rect 655 367 657 370
rect 669 369 675 375
rect 665 363 675 369
rect 710 375 720 377
rect 723 388 765 405
rect 723 387 743 388
rect 723 375 733 387
rect 738 386 741 387
rect 738 383 741 384
rect 749 384 765 388
rect 755 380 765 384
rect 751 377 752 380
rect 754 377 765 380
rect 687 367 688 370
rect 690 367 698 370
rect 700 367 702 370
rect 714 369 720 375
rect 710 363 720 369
rect 755 375 765 377
rect 768 388 810 405
rect 768 387 788 388
rect 768 375 778 387
rect 783 386 786 387
rect 783 383 786 384
rect 794 384 810 388
rect 800 380 810 384
rect 796 377 797 380
rect 799 377 810 380
rect 732 367 733 370
rect 735 367 743 370
rect 745 367 747 370
rect 759 369 765 375
rect 755 363 765 369
rect 800 375 810 377
rect 813 388 855 405
rect 813 387 833 388
rect 813 375 823 387
rect 828 386 831 387
rect 828 383 831 384
rect 839 384 855 388
rect 845 380 855 384
rect 841 377 842 380
rect 844 377 855 380
rect 777 367 778 370
rect 780 367 788 370
rect 790 367 792 370
rect 804 369 810 375
rect 800 363 810 369
rect 845 375 855 377
rect 858 388 900 405
rect 858 387 878 388
rect 858 375 868 387
rect 873 386 876 387
rect 873 383 876 384
rect 884 384 900 388
rect 890 380 900 384
rect 886 377 887 380
rect 889 377 900 380
rect 822 367 823 370
rect 825 367 833 370
rect 835 367 837 370
rect 849 369 855 375
rect 845 363 855 369
rect 890 375 900 377
rect 867 367 868 370
rect 870 367 878 370
rect 880 367 882 370
rect 894 369 900 375
rect 890 363 900 369
rect 3 343 45 360
rect 3 342 23 343
rect 3 330 13 342
rect 18 341 21 342
rect 18 338 21 339
rect 29 339 45 343
rect 35 335 45 339
rect 31 332 32 335
rect 34 332 45 335
rect 35 330 45 332
rect 48 343 90 360
rect 48 342 68 343
rect 48 330 58 342
rect 63 341 66 342
rect 63 338 66 339
rect 74 339 90 343
rect 80 335 90 339
rect 76 332 77 335
rect 79 332 90 335
rect 12 322 13 325
rect 15 322 23 325
rect 25 322 27 325
rect 39 324 45 330
rect 35 318 45 324
rect 80 330 90 332
rect 93 343 135 360
rect 93 342 113 343
rect 93 330 103 342
rect 108 341 111 342
rect 108 338 111 339
rect 119 339 135 343
rect 125 335 135 339
rect 121 332 122 335
rect 124 332 135 335
rect 57 322 58 325
rect 60 322 68 325
rect 70 322 72 325
rect 84 324 90 330
rect 80 318 90 324
rect 125 330 135 332
rect 138 343 180 360
rect 138 342 158 343
rect 138 330 148 342
rect 153 341 156 342
rect 153 338 156 339
rect 164 339 180 343
rect 170 335 180 339
rect 166 332 167 335
rect 169 332 180 335
rect 102 322 103 325
rect 105 322 113 325
rect 115 322 117 325
rect 129 324 135 330
rect 125 318 135 324
rect 170 330 180 332
rect 183 343 225 360
rect 183 342 203 343
rect 183 330 193 342
rect 198 341 201 342
rect 198 338 201 339
rect 209 339 225 343
rect 215 335 225 339
rect 211 332 212 335
rect 214 332 225 335
rect 147 322 148 325
rect 150 322 158 325
rect 160 322 162 325
rect 174 324 180 330
rect 170 318 180 324
rect 215 330 225 332
rect 228 343 270 360
rect 228 342 248 343
rect 228 330 238 342
rect 243 341 246 342
rect 243 338 246 339
rect 254 339 270 343
rect 260 335 270 339
rect 256 332 257 335
rect 259 332 270 335
rect 192 322 193 325
rect 195 322 203 325
rect 205 322 207 325
rect 219 324 225 330
rect 215 318 225 324
rect 260 330 270 332
rect 273 343 315 360
rect 273 342 293 343
rect 273 330 283 342
rect 288 341 291 342
rect 288 338 291 339
rect 299 339 315 343
rect 305 335 315 339
rect 301 332 302 335
rect 304 332 315 335
rect 237 322 238 325
rect 240 322 248 325
rect 250 322 252 325
rect 264 324 270 330
rect 260 318 270 324
rect 305 330 315 332
rect 318 343 360 360
rect 318 342 338 343
rect 318 330 328 342
rect 333 341 336 342
rect 333 338 336 339
rect 344 339 360 343
rect 350 335 360 339
rect 346 332 347 335
rect 349 332 360 335
rect 282 322 283 325
rect 285 322 293 325
rect 295 322 297 325
rect 309 324 315 330
rect 305 318 315 324
rect 350 330 360 332
rect 363 343 405 360
rect 363 342 383 343
rect 363 330 373 342
rect 378 341 381 342
rect 378 338 381 339
rect 389 339 405 343
rect 395 335 405 339
rect 391 332 392 335
rect 394 332 405 335
rect 327 322 328 325
rect 330 322 338 325
rect 340 322 342 325
rect 354 324 360 330
rect 350 318 360 324
rect 395 330 405 332
rect 408 343 450 360
rect 408 342 428 343
rect 408 330 418 342
rect 423 341 426 342
rect 423 338 426 339
rect 434 339 450 343
rect 440 335 450 339
rect 436 332 437 335
rect 439 332 450 335
rect 372 322 373 325
rect 375 322 383 325
rect 385 322 387 325
rect 399 324 405 330
rect 395 318 405 324
rect 440 330 450 332
rect 453 343 495 360
rect 453 342 473 343
rect 453 330 463 342
rect 468 341 471 342
rect 468 338 471 339
rect 479 339 495 343
rect 485 335 495 339
rect 481 332 482 335
rect 484 332 495 335
rect 417 322 418 325
rect 420 322 428 325
rect 430 322 432 325
rect 444 324 450 330
rect 440 318 450 324
rect 485 330 495 332
rect 498 343 540 360
rect 498 342 518 343
rect 498 330 508 342
rect 513 341 516 342
rect 513 338 516 339
rect 524 339 540 343
rect 530 335 540 339
rect 526 332 527 335
rect 529 332 540 335
rect 462 322 463 325
rect 465 322 473 325
rect 475 322 477 325
rect 489 324 495 330
rect 485 318 495 324
rect 530 330 540 332
rect 543 343 585 360
rect 543 342 563 343
rect 543 330 553 342
rect 558 341 561 342
rect 558 338 561 339
rect 569 339 585 343
rect 575 335 585 339
rect 571 332 572 335
rect 574 332 585 335
rect 507 322 508 325
rect 510 322 518 325
rect 520 322 522 325
rect 534 324 540 330
rect 530 318 540 324
rect 575 330 585 332
rect 588 343 630 360
rect 588 342 608 343
rect 588 330 598 342
rect 603 341 606 342
rect 603 338 606 339
rect 614 339 630 343
rect 620 335 630 339
rect 616 332 617 335
rect 619 332 630 335
rect 552 322 553 325
rect 555 322 563 325
rect 565 322 567 325
rect 579 324 585 330
rect 575 318 585 324
rect 620 330 630 332
rect 633 343 675 360
rect 633 342 653 343
rect 633 330 643 342
rect 648 341 651 342
rect 648 338 651 339
rect 659 339 675 343
rect 665 335 675 339
rect 661 332 662 335
rect 664 332 675 335
rect 597 322 598 325
rect 600 322 608 325
rect 610 322 612 325
rect 624 324 630 330
rect 620 318 630 324
rect 665 330 675 332
rect 678 343 720 360
rect 678 342 698 343
rect 678 330 688 342
rect 693 341 696 342
rect 693 338 696 339
rect 704 339 720 343
rect 710 335 720 339
rect 706 332 707 335
rect 709 332 720 335
rect 642 322 643 325
rect 645 322 653 325
rect 655 322 657 325
rect 669 324 675 330
rect 665 318 675 324
rect 710 330 720 332
rect 723 343 765 360
rect 723 342 743 343
rect 723 330 733 342
rect 738 341 741 342
rect 738 338 741 339
rect 749 339 765 343
rect 755 335 765 339
rect 751 332 752 335
rect 754 332 765 335
rect 687 322 688 325
rect 690 322 698 325
rect 700 322 702 325
rect 714 324 720 330
rect 710 318 720 324
rect 755 330 765 332
rect 768 343 810 360
rect 768 342 788 343
rect 768 330 778 342
rect 783 341 786 342
rect 783 338 786 339
rect 794 339 810 343
rect 800 335 810 339
rect 796 332 797 335
rect 799 332 810 335
rect 732 322 733 325
rect 735 322 743 325
rect 745 322 747 325
rect 759 324 765 330
rect 755 318 765 324
rect 800 330 810 332
rect 813 343 855 360
rect 813 342 833 343
rect 813 330 823 342
rect 828 341 831 342
rect 828 338 831 339
rect 839 339 855 343
rect 845 335 855 339
rect 841 332 842 335
rect 844 332 855 335
rect 777 322 778 325
rect 780 322 788 325
rect 790 322 792 325
rect 804 324 810 330
rect 800 318 810 324
rect 845 330 855 332
rect 858 343 900 360
rect 858 342 878 343
rect 858 330 868 342
rect 873 341 876 342
rect 873 338 876 339
rect 884 339 900 343
rect 890 335 900 339
rect 886 332 887 335
rect 889 332 900 335
rect 822 322 823 325
rect 825 322 833 325
rect 835 322 837 325
rect 849 324 855 330
rect 845 318 855 324
rect 890 330 900 332
rect 867 322 868 325
rect 870 322 878 325
rect 880 322 882 325
rect 894 324 900 330
rect 890 318 900 324
rect 3 298 45 315
rect 3 297 23 298
rect 3 285 13 297
rect 18 296 21 297
rect 18 293 21 294
rect 29 294 45 298
rect 35 290 45 294
rect 31 287 32 290
rect 34 287 45 290
rect 35 285 45 287
rect 48 298 90 315
rect 48 297 68 298
rect 48 285 58 297
rect 63 296 66 297
rect 63 293 66 294
rect 74 294 90 298
rect 80 290 90 294
rect 76 287 77 290
rect 79 287 90 290
rect 12 277 13 280
rect 15 277 23 280
rect 25 277 27 280
rect 39 279 45 285
rect 35 273 45 279
rect 80 285 90 287
rect 93 298 135 315
rect 93 297 113 298
rect 93 285 103 297
rect 108 296 111 297
rect 108 293 111 294
rect 119 294 135 298
rect 125 290 135 294
rect 121 287 122 290
rect 124 287 135 290
rect 57 277 58 280
rect 60 277 68 280
rect 70 277 72 280
rect 84 279 90 285
rect 80 273 90 279
rect 125 285 135 287
rect 138 298 180 315
rect 138 297 158 298
rect 138 285 148 297
rect 153 296 156 297
rect 153 293 156 294
rect 164 294 180 298
rect 170 290 180 294
rect 166 287 167 290
rect 169 287 180 290
rect 102 277 103 280
rect 105 277 113 280
rect 115 277 117 280
rect 129 279 135 285
rect 125 273 135 279
rect 170 285 180 287
rect 183 298 225 315
rect 183 297 203 298
rect 183 285 193 297
rect 198 296 201 297
rect 198 293 201 294
rect 209 294 225 298
rect 215 290 225 294
rect 211 287 212 290
rect 214 287 225 290
rect 147 277 148 280
rect 150 277 158 280
rect 160 277 162 280
rect 174 279 180 285
rect 170 273 180 279
rect 215 285 225 287
rect 228 298 270 315
rect 228 297 248 298
rect 228 285 238 297
rect 243 296 246 297
rect 243 293 246 294
rect 254 294 270 298
rect 260 290 270 294
rect 256 287 257 290
rect 259 287 270 290
rect 192 277 193 280
rect 195 277 203 280
rect 205 277 207 280
rect 219 279 225 285
rect 215 273 225 279
rect 260 285 270 287
rect 273 298 315 315
rect 273 297 293 298
rect 273 285 283 297
rect 288 296 291 297
rect 288 293 291 294
rect 299 294 315 298
rect 305 290 315 294
rect 301 287 302 290
rect 304 287 315 290
rect 237 277 238 280
rect 240 277 248 280
rect 250 277 252 280
rect 264 279 270 285
rect 260 273 270 279
rect 305 285 315 287
rect 318 298 360 315
rect 318 297 338 298
rect 318 285 328 297
rect 333 296 336 297
rect 333 293 336 294
rect 344 294 360 298
rect 350 290 360 294
rect 346 287 347 290
rect 349 287 360 290
rect 282 277 283 280
rect 285 277 293 280
rect 295 277 297 280
rect 309 279 315 285
rect 305 273 315 279
rect 350 285 360 287
rect 363 298 405 315
rect 363 297 383 298
rect 363 285 373 297
rect 378 296 381 297
rect 378 293 381 294
rect 389 294 405 298
rect 395 290 405 294
rect 391 287 392 290
rect 394 287 405 290
rect 327 277 328 280
rect 330 277 338 280
rect 340 277 342 280
rect 354 279 360 285
rect 350 273 360 279
rect 395 285 405 287
rect 408 298 450 315
rect 408 297 428 298
rect 408 285 418 297
rect 423 296 426 297
rect 423 293 426 294
rect 434 294 450 298
rect 440 290 450 294
rect 436 287 437 290
rect 439 287 450 290
rect 372 277 373 280
rect 375 277 383 280
rect 385 277 387 280
rect 399 279 405 285
rect 395 273 405 279
rect 440 285 450 287
rect 453 298 495 315
rect 453 297 473 298
rect 453 285 463 297
rect 468 296 471 297
rect 468 293 471 294
rect 479 294 495 298
rect 485 290 495 294
rect 481 287 482 290
rect 484 287 495 290
rect 417 277 418 280
rect 420 277 428 280
rect 430 277 432 280
rect 444 279 450 285
rect 440 273 450 279
rect 485 285 495 287
rect 498 298 540 315
rect 498 297 518 298
rect 498 285 508 297
rect 513 296 516 297
rect 513 293 516 294
rect 524 294 540 298
rect 530 290 540 294
rect 526 287 527 290
rect 529 287 540 290
rect 462 277 463 280
rect 465 277 473 280
rect 475 277 477 280
rect 489 279 495 285
rect 485 273 495 279
rect 530 285 540 287
rect 543 298 585 315
rect 543 297 563 298
rect 543 285 553 297
rect 558 296 561 297
rect 558 293 561 294
rect 569 294 585 298
rect 575 290 585 294
rect 571 287 572 290
rect 574 287 585 290
rect 507 277 508 280
rect 510 277 518 280
rect 520 277 522 280
rect 534 279 540 285
rect 530 273 540 279
rect 575 285 585 287
rect 588 298 630 315
rect 588 297 608 298
rect 588 285 598 297
rect 603 296 606 297
rect 603 293 606 294
rect 614 294 630 298
rect 620 290 630 294
rect 616 287 617 290
rect 619 287 630 290
rect 552 277 553 280
rect 555 277 563 280
rect 565 277 567 280
rect 579 279 585 285
rect 575 273 585 279
rect 620 285 630 287
rect 633 298 675 315
rect 633 297 653 298
rect 633 285 643 297
rect 648 296 651 297
rect 648 293 651 294
rect 659 294 675 298
rect 665 290 675 294
rect 661 287 662 290
rect 664 287 675 290
rect 597 277 598 280
rect 600 277 608 280
rect 610 277 612 280
rect 624 279 630 285
rect 620 273 630 279
rect 665 285 675 287
rect 678 298 720 315
rect 678 297 698 298
rect 678 285 688 297
rect 693 296 696 297
rect 693 293 696 294
rect 704 294 720 298
rect 710 290 720 294
rect 706 287 707 290
rect 709 287 720 290
rect 642 277 643 280
rect 645 277 653 280
rect 655 277 657 280
rect 669 279 675 285
rect 665 273 675 279
rect 710 285 720 287
rect 723 298 765 315
rect 723 297 743 298
rect 723 285 733 297
rect 738 296 741 297
rect 738 293 741 294
rect 749 294 765 298
rect 755 290 765 294
rect 751 287 752 290
rect 754 287 765 290
rect 687 277 688 280
rect 690 277 698 280
rect 700 277 702 280
rect 714 279 720 285
rect 710 273 720 279
rect 755 285 765 287
rect 768 298 810 315
rect 768 297 788 298
rect 768 285 778 297
rect 783 296 786 297
rect 783 293 786 294
rect 794 294 810 298
rect 800 290 810 294
rect 796 287 797 290
rect 799 287 810 290
rect 732 277 733 280
rect 735 277 743 280
rect 745 277 747 280
rect 759 279 765 285
rect 755 273 765 279
rect 800 285 810 287
rect 813 298 855 315
rect 813 297 833 298
rect 813 285 823 297
rect 828 296 831 297
rect 828 293 831 294
rect 839 294 855 298
rect 845 290 855 294
rect 841 287 842 290
rect 844 287 855 290
rect 777 277 778 280
rect 780 277 788 280
rect 790 277 792 280
rect 804 279 810 285
rect 800 273 810 279
rect 845 285 855 287
rect 858 298 900 315
rect 858 297 878 298
rect 858 285 868 297
rect 873 296 876 297
rect 873 293 876 294
rect 884 294 900 298
rect 890 290 900 294
rect 886 287 887 290
rect 889 287 900 290
rect 822 277 823 280
rect 825 277 833 280
rect 835 277 837 280
rect 849 279 855 285
rect 845 273 855 279
rect 890 285 900 287
rect 867 277 868 280
rect 870 277 878 280
rect 880 277 882 280
rect 894 279 900 285
rect 890 273 900 279
rect 3 253 45 270
rect 3 252 23 253
rect 3 240 13 252
rect 18 251 21 252
rect 18 248 21 249
rect 29 249 45 253
rect 35 245 45 249
rect 31 242 32 245
rect 34 242 45 245
rect 35 240 45 242
rect 48 253 90 270
rect 48 252 68 253
rect 48 240 58 252
rect 63 251 66 252
rect 63 248 66 249
rect 74 249 90 253
rect 80 245 90 249
rect 76 242 77 245
rect 79 242 90 245
rect 12 232 13 235
rect 15 232 23 235
rect 25 232 27 235
rect 39 234 45 240
rect 35 228 45 234
rect 80 240 90 242
rect 93 253 135 270
rect 93 252 113 253
rect 93 240 103 252
rect 108 251 111 252
rect 108 248 111 249
rect 119 249 135 253
rect 125 245 135 249
rect 121 242 122 245
rect 124 242 135 245
rect 57 232 58 235
rect 60 232 68 235
rect 70 232 72 235
rect 84 234 90 240
rect 80 228 90 234
rect 125 240 135 242
rect 138 253 180 270
rect 138 252 158 253
rect 138 240 148 252
rect 153 251 156 252
rect 153 248 156 249
rect 164 249 180 253
rect 170 245 180 249
rect 166 242 167 245
rect 169 242 180 245
rect 102 232 103 235
rect 105 232 113 235
rect 115 232 117 235
rect 129 234 135 240
rect 125 228 135 234
rect 170 240 180 242
rect 183 253 225 270
rect 183 252 203 253
rect 183 240 193 252
rect 198 251 201 252
rect 198 248 201 249
rect 209 249 225 253
rect 215 245 225 249
rect 211 242 212 245
rect 214 242 225 245
rect 147 232 148 235
rect 150 232 158 235
rect 160 232 162 235
rect 174 234 180 240
rect 170 228 180 234
rect 215 240 225 242
rect 228 253 270 270
rect 228 252 248 253
rect 228 240 238 252
rect 243 251 246 252
rect 243 248 246 249
rect 254 249 270 253
rect 260 245 270 249
rect 256 242 257 245
rect 259 242 270 245
rect 192 232 193 235
rect 195 232 203 235
rect 205 232 207 235
rect 219 234 225 240
rect 215 228 225 234
rect 260 240 270 242
rect 273 253 315 270
rect 273 252 293 253
rect 273 240 283 252
rect 288 251 291 252
rect 288 248 291 249
rect 299 249 315 253
rect 305 245 315 249
rect 301 242 302 245
rect 304 242 315 245
rect 237 232 238 235
rect 240 232 248 235
rect 250 232 252 235
rect 264 234 270 240
rect 260 228 270 234
rect 305 240 315 242
rect 318 253 360 270
rect 318 252 338 253
rect 318 240 328 252
rect 333 251 336 252
rect 333 248 336 249
rect 344 249 360 253
rect 350 245 360 249
rect 346 242 347 245
rect 349 242 360 245
rect 282 232 283 235
rect 285 232 293 235
rect 295 232 297 235
rect 309 234 315 240
rect 305 228 315 234
rect 350 240 360 242
rect 363 253 405 270
rect 363 252 383 253
rect 363 240 373 252
rect 378 251 381 252
rect 378 248 381 249
rect 389 249 405 253
rect 395 245 405 249
rect 391 242 392 245
rect 394 242 405 245
rect 327 232 328 235
rect 330 232 338 235
rect 340 232 342 235
rect 354 234 360 240
rect 350 228 360 234
rect 395 240 405 242
rect 408 253 450 270
rect 408 252 428 253
rect 408 240 418 252
rect 423 251 426 252
rect 423 248 426 249
rect 434 249 450 253
rect 440 245 450 249
rect 436 242 437 245
rect 439 242 450 245
rect 372 232 373 235
rect 375 232 383 235
rect 385 232 387 235
rect 399 234 405 240
rect 395 228 405 234
rect 440 240 450 242
rect 453 253 495 270
rect 453 252 473 253
rect 453 240 463 252
rect 468 251 471 252
rect 468 248 471 249
rect 479 249 495 253
rect 485 245 495 249
rect 481 242 482 245
rect 484 242 495 245
rect 417 232 418 235
rect 420 232 428 235
rect 430 232 432 235
rect 444 234 450 240
rect 440 228 450 234
rect 485 240 495 242
rect 498 253 540 270
rect 498 252 518 253
rect 498 240 508 252
rect 513 251 516 252
rect 513 248 516 249
rect 524 249 540 253
rect 530 245 540 249
rect 526 242 527 245
rect 529 242 540 245
rect 462 232 463 235
rect 465 232 473 235
rect 475 232 477 235
rect 489 234 495 240
rect 485 228 495 234
rect 530 240 540 242
rect 543 253 585 270
rect 543 252 563 253
rect 543 240 553 252
rect 558 251 561 252
rect 558 248 561 249
rect 569 249 585 253
rect 575 245 585 249
rect 571 242 572 245
rect 574 242 585 245
rect 507 232 508 235
rect 510 232 518 235
rect 520 232 522 235
rect 534 234 540 240
rect 530 228 540 234
rect 575 240 585 242
rect 588 253 630 270
rect 588 252 608 253
rect 588 240 598 252
rect 603 251 606 252
rect 603 248 606 249
rect 614 249 630 253
rect 620 245 630 249
rect 616 242 617 245
rect 619 242 630 245
rect 552 232 553 235
rect 555 232 563 235
rect 565 232 567 235
rect 579 234 585 240
rect 575 228 585 234
rect 620 240 630 242
rect 633 253 675 270
rect 633 252 653 253
rect 633 240 643 252
rect 648 251 651 252
rect 648 248 651 249
rect 659 249 675 253
rect 665 245 675 249
rect 661 242 662 245
rect 664 242 675 245
rect 597 232 598 235
rect 600 232 608 235
rect 610 232 612 235
rect 624 234 630 240
rect 620 228 630 234
rect 665 240 675 242
rect 678 253 720 270
rect 678 252 698 253
rect 678 240 688 252
rect 693 251 696 252
rect 693 248 696 249
rect 704 249 720 253
rect 710 245 720 249
rect 706 242 707 245
rect 709 242 720 245
rect 642 232 643 235
rect 645 232 653 235
rect 655 232 657 235
rect 669 234 675 240
rect 665 228 675 234
rect 710 240 720 242
rect 723 253 765 270
rect 723 252 743 253
rect 723 240 733 252
rect 738 251 741 252
rect 738 248 741 249
rect 749 249 765 253
rect 755 245 765 249
rect 751 242 752 245
rect 754 242 765 245
rect 687 232 688 235
rect 690 232 698 235
rect 700 232 702 235
rect 714 234 720 240
rect 710 228 720 234
rect 755 240 765 242
rect 768 253 810 270
rect 768 252 788 253
rect 768 240 778 252
rect 783 251 786 252
rect 783 248 786 249
rect 794 249 810 253
rect 800 245 810 249
rect 796 242 797 245
rect 799 242 810 245
rect 732 232 733 235
rect 735 232 743 235
rect 745 232 747 235
rect 759 234 765 240
rect 755 228 765 234
rect 800 240 810 242
rect 813 253 855 270
rect 813 252 833 253
rect 813 240 823 252
rect 828 251 831 252
rect 828 248 831 249
rect 839 249 855 253
rect 845 245 855 249
rect 841 242 842 245
rect 844 242 855 245
rect 777 232 778 235
rect 780 232 788 235
rect 790 232 792 235
rect 804 234 810 240
rect 800 228 810 234
rect 845 240 855 242
rect 858 253 900 270
rect 858 252 878 253
rect 858 240 868 252
rect 873 251 876 252
rect 873 248 876 249
rect 884 249 900 253
rect 890 245 900 249
rect 886 242 887 245
rect 889 242 900 245
rect 822 232 823 235
rect 825 232 833 235
rect 835 232 837 235
rect 849 234 855 240
rect 845 228 855 234
rect 890 240 900 242
rect 867 232 868 235
rect 870 232 878 235
rect 880 232 882 235
rect 894 234 900 240
rect 890 228 900 234
rect 3 208 45 225
rect 3 207 23 208
rect 3 195 13 207
rect 18 206 21 207
rect 18 203 21 204
rect 29 204 45 208
rect 35 200 45 204
rect 31 197 32 200
rect 34 197 45 200
rect 35 195 45 197
rect 48 208 90 225
rect 48 207 68 208
rect 48 195 58 207
rect 63 206 66 207
rect 63 203 66 204
rect 74 204 90 208
rect 80 200 90 204
rect 76 197 77 200
rect 79 197 90 200
rect 12 187 13 190
rect 15 187 23 190
rect 25 187 27 190
rect 39 189 45 195
rect 35 183 45 189
rect 80 195 90 197
rect 93 208 135 225
rect 93 207 113 208
rect 93 195 103 207
rect 108 206 111 207
rect 108 203 111 204
rect 119 204 135 208
rect 125 200 135 204
rect 121 197 122 200
rect 124 197 135 200
rect 57 187 58 190
rect 60 187 68 190
rect 70 187 72 190
rect 84 189 90 195
rect 80 183 90 189
rect 125 195 135 197
rect 138 208 180 225
rect 138 207 158 208
rect 138 195 148 207
rect 153 206 156 207
rect 153 203 156 204
rect 164 204 180 208
rect 170 200 180 204
rect 166 197 167 200
rect 169 197 180 200
rect 102 187 103 190
rect 105 187 113 190
rect 115 187 117 190
rect 129 189 135 195
rect 125 183 135 189
rect 170 195 180 197
rect 183 208 225 225
rect 183 207 203 208
rect 183 195 193 207
rect 198 206 201 207
rect 198 203 201 204
rect 209 204 225 208
rect 215 200 225 204
rect 211 197 212 200
rect 214 197 225 200
rect 147 187 148 190
rect 150 187 158 190
rect 160 187 162 190
rect 174 189 180 195
rect 170 183 180 189
rect 215 195 225 197
rect 228 208 270 225
rect 228 207 248 208
rect 228 195 238 207
rect 243 206 246 207
rect 243 203 246 204
rect 254 204 270 208
rect 260 200 270 204
rect 256 197 257 200
rect 259 197 270 200
rect 192 187 193 190
rect 195 187 203 190
rect 205 187 207 190
rect 219 189 225 195
rect 215 183 225 189
rect 260 195 270 197
rect 273 208 315 225
rect 273 207 293 208
rect 273 195 283 207
rect 288 206 291 207
rect 288 203 291 204
rect 299 204 315 208
rect 305 200 315 204
rect 301 197 302 200
rect 304 197 315 200
rect 237 187 238 190
rect 240 187 248 190
rect 250 187 252 190
rect 264 189 270 195
rect 260 183 270 189
rect 305 195 315 197
rect 318 208 360 225
rect 318 207 338 208
rect 318 195 328 207
rect 333 206 336 207
rect 333 203 336 204
rect 344 204 360 208
rect 350 200 360 204
rect 346 197 347 200
rect 349 197 360 200
rect 282 187 283 190
rect 285 187 293 190
rect 295 187 297 190
rect 309 189 315 195
rect 305 183 315 189
rect 350 195 360 197
rect 363 208 405 225
rect 363 207 383 208
rect 363 195 373 207
rect 378 206 381 207
rect 378 203 381 204
rect 389 204 405 208
rect 395 200 405 204
rect 391 197 392 200
rect 394 197 405 200
rect 327 187 328 190
rect 330 187 338 190
rect 340 187 342 190
rect 354 189 360 195
rect 350 183 360 189
rect 395 195 405 197
rect 408 208 450 225
rect 408 207 428 208
rect 408 195 418 207
rect 423 206 426 207
rect 423 203 426 204
rect 434 204 450 208
rect 440 200 450 204
rect 436 197 437 200
rect 439 197 450 200
rect 372 187 373 190
rect 375 187 383 190
rect 385 187 387 190
rect 399 189 405 195
rect 395 183 405 189
rect 440 195 450 197
rect 453 208 495 225
rect 453 207 473 208
rect 453 195 463 207
rect 468 206 471 207
rect 468 203 471 204
rect 479 204 495 208
rect 485 200 495 204
rect 481 197 482 200
rect 484 197 495 200
rect 417 187 418 190
rect 420 187 428 190
rect 430 187 432 190
rect 444 189 450 195
rect 440 183 450 189
rect 485 195 495 197
rect 498 208 540 225
rect 498 207 518 208
rect 498 195 508 207
rect 513 206 516 207
rect 513 203 516 204
rect 524 204 540 208
rect 530 200 540 204
rect 526 197 527 200
rect 529 197 540 200
rect 462 187 463 190
rect 465 187 473 190
rect 475 187 477 190
rect 489 189 495 195
rect 485 183 495 189
rect 530 195 540 197
rect 543 208 585 225
rect 543 207 563 208
rect 543 195 553 207
rect 558 206 561 207
rect 558 203 561 204
rect 569 204 585 208
rect 575 200 585 204
rect 571 197 572 200
rect 574 197 585 200
rect 507 187 508 190
rect 510 187 518 190
rect 520 187 522 190
rect 534 189 540 195
rect 530 183 540 189
rect 575 195 585 197
rect 588 208 630 225
rect 588 207 608 208
rect 588 195 598 207
rect 603 206 606 207
rect 603 203 606 204
rect 614 204 630 208
rect 620 200 630 204
rect 616 197 617 200
rect 619 197 630 200
rect 552 187 553 190
rect 555 187 563 190
rect 565 187 567 190
rect 579 189 585 195
rect 575 183 585 189
rect 620 195 630 197
rect 633 208 675 225
rect 633 207 653 208
rect 633 195 643 207
rect 648 206 651 207
rect 648 203 651 204
rect 659 204 675 208
rect 665 200 675 204
rect 661 197 662 200
rect 664 197 675 200
rect 597 187 598 190
rect 600 187 608 190
rect 610 187 612 190
rect 624 189 630 195
rect 620 183 630 189
rect 665 195 675 197
rect 678 208 720 225
rect 678 207 698 208
rect 678 195 688 207
rect 693 206 696 207
rect 693 203 696 204
rect 704 204 720 208
rect 710 200 720 204
rect 706 197 707 200
rect 709 197 720 200
rect 642 187 643 190
rect 645 187 653 190
rect 655 187 657 190
rect 669 189 675 195
rect 665 183 675 189
rect 710 195 720 197
rect 723 208 765 225
rect 723 207 743 208
rect 723 195 733 207
rect 738 206 741 207
rect 738 203 741 204
rect 749 204 765 208
rect 755 200 765 204
rect 751 197 752 200
rect 754 197 765 200
rect 687 187 688 190
rect 690 187 698 190
rect 700 187 702 190
rect 714 189 720 195
rect 710 183 720 189
rect 755 195 765 197
rect 768 208 810 225
rect 768 207 788 208
rect 768 195 778 207
rect 783 206 786 207
rect 783 203 786 204
rect 794 204 810 208
rect 800 200 810 204
rect 796 197 797 200
rect 799 197 810 200
rect 732 187 733 190
rect 735 187 743 190
rect 745 187 747 190
rect 759 189 765 195
rect 755 183 765 189
rect 800 195 810 197
rect 813 208 855 225
rect 813 207 833 208
rect 813 195 823 207
rect 828 206 831 207
rect 828 203 831 204
rect 839 204 855 208
rect 845 200 855 204
rect 841 197 842 200
rect 844 197 855 200
rect 777 187 778 190
rect 780 187 788 190
rect 790 187 792 190
rect 804 189 810 195
rect 800 183 810 189
rect 845 195 855 197
rect 858 208 900 225
rect 858 207 878 208
rect 858 195 868 207
rect 873 206 876 207
rect 873 203 876 204
rect 884 204 900 208
rect 890 200 900 204
rect 886 197 887 200
rect 889 197 900 200
rect 822 187 823 190
rect 825 187 833 190
rect 835 187 837 190
rect 849 189 855 195
rect 845 183 855 189
rect 890 195 900 197
rect 867 187 868 190
rect 870 187 878 190
rect 880 187 882 190
rect 894 189 900 195
rect 890 183 900 189
rect 3 163 45 180
rect 3 162 23 163
rect 3 150 13 162
rect 18 161 21 162
rect 18 158 21 159
rect 29 159 45 163
rect 35 155 45 159
rect 31 152 32 155
rect 34 152 45 155
rect 35 150 45 152
rect 48 163 90 180
rect 48 162 68 163
rect 48 150 58 162
rect 63 161 66 162
rect 63 158 66 159
rect 74 159 90 163
rect 80 155 90 159
rect 76 152 77 155
rect 79 152 90 155
rect 12 142 13 145
rect 15 142 23 145
rect 25 142 27 145
rect 39 144 45 150
rect 35 138 45 144
rect 80 150 90 152
rect 93 163 135 180
rect 93 162 113 163
rect 93 150 103 162
rect 108 161 111 162
rect 108 158 111 159
rect 119 159 135 163
rect 125 155 135 159
rect 121 152 122 155
rect 124 152 135 155
rect 57 142 58 145
rect 60 142 68 145
rect 70 142 72 145
rect 84 144 90 150
rect 80 138 90 144
rect 125 150 135 152
rect 138 163 180 180
rect 138 162 158 163
rect 138 150 148 162
rect 153 161 156 162
rect 153 158 156 159
rect 164 159 180 163
rect 170 155 180 159
rect 166 152 167 155
rect 169 152 180 155
rect 102 142 103 145
rect 105 142 113 145
rect 115 142 117 145
rect 129 144 135 150
rect 125 138 135 144
rect 170 150 180 152
rect 183 163 225 180
rect 183 162 203 163
rect 183 150 193 162
rect 198 161 201 162
rect 198 158 201 159
rect 209 159 225 163
rect 215 155 225 159
rect 211 152 212 155
rect 214 152 225 155
rect 147 142 148 145
rect 150 142 158 145
rect 160 142 162 145
rect 174 144 180 150
rect 170 138 180 144
rect 215 150 225 152
rect 228 163 270 180
rect 228 162 248 163
rect 228 150 238 162
rect 243 161 246 162
rect 243 158 246 159
rect 254 159 270 163
rect 260 155 270 159
rect 256 152 257 155
rect 259 152 270 155
rect 192 142 193 145
rect 195 142 203 145
rect 205 142 207 145
rect 219 144 225 150
rect 215 138 225 144
rect 260 150 270 152
rect 273 163 315 180
rect 273 162 293 163
rect 273 150 283 162
rect 288 161 291 162
rect 288 158 291 159
rect 299 159 315 163
rect 305 155 315 159
rect 301 152 302 155
rect 304 152 315 155
rect 237 142 238 145
rect 240 142 248 145
rect 250 142 252 145
rect 264 144 270 150
rect 260 138 270 144
rect 305 150 315 152
rect 318 163 360 180
rect 318 162 338 163
rect 318 150 328 162
rect 333 161 336 162
rect 333 158 336 159
rect 344 159 360 163
rect 350 155 360 159
rect 346 152 347 155
rect 349 152 360 155
rect 282 142 283 145
rect 285 142 293 145
rect 295 142 297 145
rect 309 144 315 150
rect 305 138 315 144
rect 350 150 360 152
rect 363 163 405 180
rect 363 162 383 163
rect 363 150 373 162
rect 378 161 381 162
rect 378 158 381 159
rect 389 159 405 163
rect 395 155 405 159
rect 391 152 392 155
rect 394 152 405 155
rect 327 142 328 145
rect 330 142 338 145
rect 340 142 342 145
rect 354 144 360 150
rect 350 138 360 144
rect 395 150 405 152
rect 408 163 450 180
rect 408 162 428 163
rect 408 150 418 162
rect 423 161 426 162
rect 423 158 426 159
rect 434 159 450 163
rect 440 155 450 159
rect 436 152 437 155
rect 439 152 450 155
rect 372 142 373 145
rect 375 142 383 145
rect 385 142 387 145
rect 399 144 405 150
rect 395 138 405 144
rect 440 150 450 152
rect 453 163 495 180
rect 453 162 473 163
rect 453 150 463 162
rect 468 161 471 162
rect 468 158 471 159
rect 479 159 495 163
rect 485 155 495 159
rect 481 152 482 155
rect 484 152 495 155
rect 417 142 418 145
rect 420 142 428 145
rect 430 142 432 145
rect 444 144 450 150
rect 440 138 450 144
rect 485 150 495 152
rect 498 163 540 180
rect 498 162 518 163
rect 498 150 508 162
rect 513 161 516 162
rect 513 158 516 159
rect 524 159 540 163
rect 530 155 540 159
rect 526 152 527 155
rect 529 152 540 155
rect 462 142 463 145
rect 465 142 473 145
rect 475 142 477 145
rect 489 144 495 150
rect 485 138 495 144
rect 530 150 540 152
rect 543 163 585 180
rect 543 162 563 163
rect 543 150 553 162
rect 558 161 561 162
rect 558 158 561 159
rect 569 159 585 163
rect 575 155 585 159
rect 571 152 572 155
rect 574 152 585 155
rect 507 142 508 145
rect 510 142 518 145
rect 520 142 522 145
rect 534 144 540 150
rect 530 138 540 144
rect 575 150 585 152
rect 588 163 630 180
rect 588 162 608 163
rect 588 150 598 162
rect 603 161 606 162
rect 603 158 606 159
rect 614 159 630 163
rect 620 155 630 159
rect 616 152 617 155
rect 619 152 630 155
rect 552 142 553 145
rect 555 142 563 145
rect 565 142 567 145
rect 579 144 585 150
rect 575 138 585 144
rect 620 150 630 152
rect 633 163 675 180
rect 633 162 653 163
rect 633 150 643 162
rect 648 161 651 162
rect 648 158 651 159
rect 659 159 675 163
rect 665 155 675 159
rect 661 152 662 155
rect 664 152 675 155
rect 597 142 598 145
rect 600 142 608 145
rect 610 142 612 145
rect 624 144 630 150
rect 620 138 630 144
rect 665 150 675 152
rect 678 163 720 180
rect 678 162 698 163
rect 678 150 688 162
rect 693 161 696 162
rect 693 158 696 159
rect 704 159 720 163
rect 710 155 720 159
rect 706 152 707 155
rect 709 152 720 155
rect 642 142 643 145
rect 645 142 653 145
rect 655 142 657 145
rect 669 144 675 150
rect 665 138 675 144
rect 710 150 720 152
rect 723 163 765 180
rect 723 162 743 163
rect 723 150 733 162
rect 738 161 741 162
rect 738 158 741 159
rect 749 159 765 163
rect 755 155 765 159
rect 751 152 752 155
rect 754 152 765 155
rect 687 142 688 145
rect 690 142 698 145
rect 700 142 702 145
rect 714 144 720 150
rect 710 138 720 144
rect 755 150 765 152
rect 768 163 810 180
rect 768 162 788 163
rect 768 150 778 162
rect 783 161 786 162
rect 783 158 786 159
rect 794 159 810 163
rect 800 155 810 159
rect 796 152 797 155
rect 799 152 810 155
rect 732 142 733 145
rect 735 142 743 145
rect 745 142 747 145
rect 759 144 765 150
rect 755 138 765 144
rect 800 150 810 152
rect 813 163 855 180
rect 813 162 833 163
rect 813 150 823 162
rect 828 161 831 162
rect 828 158 831 159
rect 839 159 855 163
rect 845 155 855 159
rect 841 152 842 155
rect 844 152 855 155
rect 777 142 778 145
rect 780 142 788 145
rect 790 142 792 145
rect 804 144 810 150
rect 800 138 810 144
rect 845 150 855 152
rect 858 163 900 180
rect 858 162 878 163
rect 858 150 868 162
rect 873 161 876 162
rect 873 158 876 159
rect 884 159 900 163
rect 890 155 900 159
rect 886 152 887 155
rect 889 152 900 155
rect 822 142 823 145
rect 825 142 833 145
rect 835 142 837 145
rect 849 144 855 150
rect 845 138 855 144
rect 890 150 900 152
rect 867 142 868 145
rect 870 142 878 145
rect 880 142 882 145
rect 894 144 900 150
rect 890 138 900 144
rect 3 118 45 135
rect 3 117 23 118
rect 3 105 13 117
rect 18 116 21 117
rect 18 113 21 114
rect 29 114 45 118
rect 35 110 45 114
rect 31 107 32 110
rect 34 107 45 110
rect 35 105 45 107
rect 48 118 90 135
rect 48 117 68 118
rect 48 105 58 117
rect 63 116 66 117
rect 63 113 66 114
rect 74 114 90 118
rect 80 110 90 114
rect 76 107 77 110
rect 79 107 90 110
rect 12 97 13 100
rect 15 97 23 100
rect 25 97 27 100
rect 39 99 45 105
rect 35 93 45 99
rect 80 105 90 107
rect 93 118 135 135
rect 93 117 113 118
rect 93 105 103 117
rect 108 116 111 117
rect 108 113 111 114
rect 119 114 135 118
rect 125 110 135 114
rect 121 107 122 110
rect 124 107 135 110
rect 57 97 58 100
rect 60 97 68 100
rect 70 97 72 100
rect 84 99 90 105
rect 80 93 90 99
rect 125 105 135 107
rect 138 118 180 135
rect 138 117 158 118
rect 138 105 148 117
rect 153 116 156 117
rect 153 113 156 114
rect 164 114 180 118
rect 170 110 180 114
rect 166 107 167 110
rect 169 107 180 110
rect 102 97 103 100
rect 105 97 113 100
rect 115 97 117 100
rect 129 99 135 105
rect 125 93 135 99
rect 170 105 180 107
rect 183 118 225 135
rect 183 117 203 118
rect 183 105 193 117
rect 198 116 201 117
rect 198 113 201 114
rect 209 114 225 118
rect 215 110 225 114
rect 211 107 212 110
rect 214 107 225 110
rect 147 97 148 100
rect 150 97 158 100
rect 160 97 162 100
rect 174 99 180 105
rect 170 93 180 99
rect 215 105 225 107
rect 228 118 270 135
rect 228 117 248 118
rect 228 105 238 117
rect 243 116 246 117
rect 243 113 246 114
rect 254 114 270 118
rect 260 110 270 114
rect 256 107 257 110
rect 259 107 270 110
rect 192 97 193 100
rect 195 97 203 100
rect 205 97 207 100
rect 219 99 225 105
rect 215 93 225 99
rect 260 105 270 107
rect 273 118 315 135
rect 273 117 293 118
rect 273 105 283 117
rect 288 116 291 117
rect 288 113 291 114
rect 299 114 315 118
rect 305 110 315 114
rect 301 107 302 110
rect 304 107 315 110
rect 237 97 238 100
rect 240 97 248 100
rect 250 97 252 100
rect 264 99 270 105
rect 260 93 270 99
rect 305 105 315 107
rect 318 118 360 135
rect 318 117 338 118
rect 318 105 328 117
rect 333 116 336 117
rect 333 113 336 114
rect 344 114 360 118
rect 350 110 360 114
rect 346 107 347 110
rect 349 107 360 110
rect 282 97 283 100
rect 285 97 293 100
rect 295 97 297 100
rect 309 99 315 105
rect 305 93 315 99
rect 350 105 360 107
rect 363 118 405 135
rect 363 117 383 118
rect 363 105 373 117
rect 378 116 381 117
rect 378 113 381 114
rect 389 114 405 118
rect 395 110 405 114
rect 391 107 392 110
rect 394 107 405 110
rect 327 97 328 100
rect 330 97 338 100
rect 340 97 342 100
rect 354 99 360 105
rect 350 93 360 99
rect 395 105 405 107
rect 408 118 450 135
rect 408 117 428 118
rect 408 105 418 117
rect 423 116 426 117
rect 423 113 426 114
rect 434 114 450 118
rect 440 110 450 114
rect 436 107 437 110
rect 439 107 450 110
rect 372 97 373 100
rect 375 97 383 100
rect 385 97 387 100
rect 399 99 405 105
rect 395 93 405 99
rect 440 105 450 107
rect 453 118 495 135
rect 453 117 473 118
rect 453 105 463 117
rect 468 116 471 117
rect 468 113 471 114
rect 479 114 495 118
rect 485 110 495 114
rect 481 107 482 110
rect 484 107 495 110
rect 417 97 418 100
rect 420 97 428 100
rect 430 97 432 100
rect 444 99 450 105
rect 440 93 450 99
rect 485 105 495 107
rect 498 118 540 135
rect 498 117 518 118
rect 498 105 508 117
rect 513 116 516 117
rect 513 113 516 114
rect 524 114 540 118
rect 530 110 540 114
rect 526 107 527 110
rect 529 107 540 110
rect 462 97 463 100
rect 465 97 473 100
rect 475 97 477 100
rect 489 99 495 105
rect 485 93 495 99
rect 530 105 540 107
rect 543 118 585 135
rect 543 117 563 118
rect 543 105 553 117
rect 558 116 561 117
rect 558 113 561 114
rect 569 114 585 118
rect 575 110 585 114
rect 571 107 572 110
rect 574 107 585 110
rect 507 97 508 100
rect 510 97 518 100
rect 520 97 522 100
rect 534 99 540 105
rect 530 93 540 99
rect 575 105 585 107
rect 588 118 630 135
rect 588 117 608 118
rect 588 105 598 117
rect 603 116 606 117
rect 603 113 606 114
rect 614 114 630 118
rect 620 110 630 114
rect 616 107 617 110
rect 619 107 630 110
rect 552 97 553 100
rect 555 97 563 100
rect 565 97 567 100
rect 579 99 585 105
rect 575 93 585 99
rect 620 105 630 107
rect 633 118 675 135
rect 633 117 653 118
rect 633 105 643 117
rect 648 116 651 117
rect 648 113 651 114
rect 659 114 675 118
rect 665 110 675 114
rect 661 107 662 110
rect 664 107 675 110
rect 597 97 598 100
rect 600 97 608 100
rect 610 97 612 100
rect 624 99 630 105
rect 620 93 630 99
rect 665 105 675 107
rect 678 118 720 135
rect 678 117 698 118
rect 678 105 688 117
rect 693 116 696 117
rect 693 113 696 114
rect 704 114 720 118
rect 710 110 720 114
rect 706 107 707 110
rect 709 107 720 110
rect 642 97 643 100
rect 645 97 653 100
rect 655 97 657 100
rect 669 99 675 105
rect 665 93 675 99
rect 710 105 720 107
rect 723 118 765 135
rect 723 117 743 118
rect 723 105 733 117
rect 738 116 741 117
rect 738 113 741 114
rect 749 114 765 118
rect 755 110 765 114
rect 751 107 752 110
rect 754 107 765 110
rect 687 97 688 100
rect 690 97 698 100
rect 700 97 702 100
rect 714 99 720 105
rect 710 93 720 99
rect 755 105 765 107
rect 768 118 810 135
rect 768 117 788 118
rect 768 105 778 117
rect 783 116 786 117
rect 783 113 786 114
rect 794 114 810 118
rect 800 110 810 114
rect 796 107 797 110
rect 799 107 810 110
rect 732 97 733 100
rect 735 97 743 100
rect 745 97 747 100
rect 759 99 765 105
rect 755 93 765 99
rect 800 105 810 107
rect 813 118 855 135
rect 813 117 833 118
rect 813 105 823 117
rect 828 116 831 117
rect 828 113 831 114
rect 839 114 855 118
rect 845 110 855 114
rect 841 107 842 110
rect 844 107 855 110
rect 777 97 778 100
rect 780 97 788 100
rect 790 97 792 100
rect 804 99 810 105
rect 800 93 810 99
rect 845 105 855 107
rect 858 118 900 135
rect 858 117 878 118
rect 858 105 868 117
rect 873 116 876 117
rect 873 113 876 114
rect 884 114 900 118
rect 890 110 900 114
rect 886 107 887 110
rect 889 107 900 110
rect 822 97 823 100
rect 825 97 833 100
rect 835 97 837 100
rect 849 99 855 105
rect 845 93 855 99
rect 890 105 900 107
rect 867 97 868 100
rect 870 97 878 100
rect 880 97 882 100
rect 894 99 900 105
rect 890 93 900 99
rect 3 73 45 90
rect 3 72 23 73
rect 3 60 13 72
rect 18 71 21 72
rect 18 68 21 69
rect 29 69 45 73
rect 35 65 45 69
rect 31 62 32 65
rect 34 62 45 65
rect 35 60 45 62
rect 48 73 90 90
rect 48 72 68 73
rect 48 60 58 72
rect 63 71 66 72
rect 63 68 66 69
rect 74 69 90 73
rect 80 65 90 69
rect 76 62 77 65
rect 79 62 90 65
rect 12 52 13 55
rect 15 52 23 55
rect 25 52 27 55
rect 39 54 45 60
rect 35 48 45 54
rect 80 60 90 62
rect 93 73 135 90
rect 93 72 113 73
rect 93 60 103 72
rect 108 71 111 72
rect 108 68 111 69
rect 119 69 135 73
rect 125 65 135 69
rect 121 62 122 65
rect 124 62 135 65
rect 57 52 58 55
rect 60 52 68 55
rect 70 52 72 55
rect 84 54 90 60
rect 80 48 90 54
rect 125 60 135 62
rect 138 73 180 90
rect 138 72 158 73
rect 138 60 148 72
rect 153 71 156 72
rect 153 68 156 69
rect 164 69 180 73
rect 170 65 180 69
rect 166 62 167 65
rect 169 62 180 65
rect 102 52 103 55
rect 105 52 113 55
rect 115 52 117 55
rect 129 54 135 60
rect 125 48 135 54
rect 170 60 180 62
rect 183 73 225 90
rect 183 72 203 73
rect 183 60 193 72
rect 198 71 201 72
rect 198 68 201 69
rect 209 69 225 73
rect 215 65 225 69
rect 211 62 212 65
rect 214 62 225 65
rect 147 52 148 55
rect 150 52 158 55
rect 160 52 162 55
rect 174 54 180 60
rect 170 48 180 54
rect 215 60 225 62
rect 228 73 270 90
rect 228 72 248 73
rect 228 60 238 72
rect 243 71 246 72
rect 243 68 246 69
rect 254 69 270 73
rect 260 65 270 69
rect 256 62 257 65
rect 259 62 270 65
rect 192 52 193 55
rect 195 52 203 55
rect 205 52 207 55
rect 219 54 225 60
rect 215 48 225 54
rect 260 60 270 62
rect 273 73 315 90
rect 273 72 293 73
rect 273 60 283 72
rect 288 71 291 72
rect 288 68 291 69
rect 299 69 315 73
rect 305 65 315 69
rect 301 62 302 65
rect 304 62 315 65
rect 237 52 238 55
rect 240 52 248 55
rect 250 52 252 55
rect 264 54 270 60
rect 260 48 270 54
rect 305 60 315 62
rect 318 73 360 90
rect 318 72 338 73
rect 318 60 328 72
rect 333 71 336 72
rect 333 68 336 69
rect 344 69 360 73
rect 350 65 360 69
rect 346 62 347 65
rect 349 62 360 65
rect 282 52 283 55
rect 285 52 293 55
rect 295 52 297 55
rect 309 54 315 60
rect 305 48 315 54
rect 350 60 360 62
rect 363 73 405 90
rect 363 72 383 73
rect 363 60 373 72
rect 378 71 381 72
rect 378 68 381 69
rect 389 69 405 73
rect 395 65 405 69
rect 391 62 392 65
rect 394 62 405 65
rect 327 52 328 55
rect 330 52 338 55
rect 340 52 342 55
rect 354 54 360 60
rect 350 48 360 54
rect 395 60 405 62
rect 408 73 450 90
rect 408 72 428 73
rect 408 60 418 72
rect 423 71 426 72
rect 423 68 426 69
rect 434 69 450 73
rect 440 65 450 69
rect 436 62 437 65
rect 439 62 450 65
rect 372 52 373 55
rect 375 52 383 55
rect 385 52 387 55
rect 399 54 405 60
rect 395 48 405 54
rect 440 60 450 62
rect 453 73 495 90
rect 453 72 473 73
rect 453 60 463 72
rect 468 71 471 72
rect 468 68 471 69
rect 479 69 495 73
rect 485 65 495 69
rect 481 62 482 65
rect 484 62 495 65
rect 417 52 418 55
rect 420 52 428 55
rect 430 52 432 55
rect 444 54 450 60
rect 440 48 450 54
rect 485 60 495 62
rect 498 73 540 90
rect 498 72 518 73
rect 498 60 508 72
rect 513 71 516 72
rect 513 68 516 69
rect 524 69 540 73
rect 530 65 540 69
rect 526 62 527 65
rect 529 62 540 65
rect 462 52 463 55
rect 465 52 473 55
rect 475 52 477 55
rect 489 54 495 60
rect 485 48 495 54
rect 530 60 540 62
rect 543 73 585 90
rect 543 72 563 73
rect 543 60 553 72
rect 558 71 561 72
rect 558 68 561 69
rect 569 69 585 73
rect 575 65 585 69
rect 571 62 572 65
rect 574 62 585 65
rect 507 52 508 55
rect 510 52 518 55
rect 520 52 522 55
rect 534 54 540 60
rect 530 48 540 54
rect 575 60 585 62
rect 588 73 630 90
rect 588 72 608 73
rect 588 60 598 72
rect 603 71 606 72
rect 603 68 606 69
rect 614 69 630 73
rect 620 65 630 69
rect 616 62 617 65
rect 619 62 630 65
rect 552 52 553 55
rect 555 52 563 55
rect 565 52 567 55
rect 579 54 585 60
rect 575 48 585 54
rect 620 60 630 62
rect 633 73 675 90
rect 633 72 653 73
rect 633 60 643 72
rect 648 71 651 72
rect 648 68 651 69
rect 659 69 675 73
rect 665 65 675 69
rect 661 62 662 65
rect 664 62 675 65
rect 597 52 598 55
rect 600 52 608 55
rect 610 52 612 55
rect 624 54 630 60
rect 620 48 630 54
rect 665 60 675 62
rect 678 73 720 90
rect 678 72 698 73
rect 678 60 688 72
rect 693 71 696 72
rect 693 68 696 69
rect 704 69 720 73
rect 710 65 720 69
rect 706 62 707 65
rect 709 62 720 65
rect 642 52 643 55
rect 645 52 653 55
rect 655 52 657 55
rect 669 54 675 60
rect 665 48 675 54
rect 710 60 720 62
rect 723 73 765 90
rect 723 72 743 73
rect 723 60 733 72
rect 738 71 741 72
rect 738 68 741 69
rect 749 69 765 73
rect 755 65 765 69
rect 751 62 752 65
rect 754 62 765 65
rect 687 52 688 55
rect 690 52 698 55
rect 700 52 702 55
rect 714 54 720 60
rect 710 48 720 54
rect 755 60 765 62
rect 768 73 810 90
rect 768 72 788 73
rect 768 60 778 72
rect 783 71 786 72
rect 783 68 786 69
rect 794 69 810 73
rect 800 65 810 69
rect 796 62 797 65
rect 799 62 810 65
rect 732 52 733 55
rect 735 52 743 55
rect 745 52 747 55
rect 759 54 765 60
rect 755 48 765 54
rect 800 60 810 62
rect 813 73 855 90
rect 813 72 833 73
rect 813 60 823 72
rect 828 71 831 72
rect 828 68 831 69
rect 839 69 855 73
rect 845 65 855 69
rect 841 62 842 65
rect 844 62 855 65
rect 777 52 778 55
rect 780 52 788 55
rect 790 52 792 55
rect 804 54 810 60
rect 800 48 810 54
rect 845 60 855 62
rect 858 73 900 90
rect 858 72 878 73
rect 858 60 868 72
rect 873 71 876 72
rect 873 68 876 69
rect 884 69 900 73
rect 890 65 900 69
rect 886 62 887 65
rect 889 62 900 65
rect 822 52 823 55
rect 825 52 833 55
rect 835 52 837 55
rect 849 54 855 60
rect 845 48 855 54
rect 890 60 900 62
rect 867 52 868 55
rect 870 52 878 55
rect 880 52 882 55
rect 894 54 900 60
rect 890 48 900 54
rect 3 28 45 45
rect 3 27 23 28
rect 3 15 13 27
rect 18 26 21 27
rect 18 23 21 24
rect 29 24 45 28
rect 35 20 45 24
rect 31 17 32 20
rect 34 17 45 20
rect 35 15 45 17
rect 48 28 90 45
rect 48 27 68 28
rect 48 15 58 27
rect 63 26 66 27
rect 63 23 66 24
rect 74 24 90 28
rect 80 20 90 24
rect 76 17 77 20
rect 79 17 90 20
rect 12 7 13 10
rect 15 7 23 10
rect 25 7 27 10
rect 39 9 45 15
rect 35 3 45 9
rect 80 15 90 17
rect 93 28 135 45
rect 93 27 113 28
rect 93 15 103 27
rect 108 26 111 27
rect 108 23 111 24
rect 119 24 135 28
rect 125 20 135 24
rect 121 17 122 20
rect 124 17 135 20
rect 57 7 58 10
rect 60 7 68 10
rect 70 7 72 10
rect 84 9 90 15
rect 80 3 90 9
rect 125 15 135 17
rect 138 28 180 45
rect 138 27 158 28
rect 138 15 148 27
rect 153 26 156 27
rect 153 23 156 24
rect 164 24 180 28
rect 170 20 180 24
rect 166 17 167 20
rect 169 17 180 20
rect 102 7 103 10
rect 105 7 113 10
rect 115 7 117 10
rect 129 9 135 15
rect 125 3 135 9
rect 170 15 180 17
rect 183 28 225 45
rect 183 27 203 28
rect 183 15 193 27
rect 198 26 201 27
rect 198 23 201 24
rect 209 24 225 28
rect 215 20 225 24
rect 211 17 212 20
rect 214 17 225 20
rect 147 7 148 10
rect 150 7 158 10
rect 160 7 162 10
rect 174 9 180 15
rect 170 3 180 9
rect 215 15 225 17
rect 228 28 270 45
rect 228 27 248 28
rect 228 15 238 27
rect 243 26 246 27
rect 243 23 246 24
rect 254 24 270 28
rect 260 20 270 24
rect 256 17 257 20
rect 259 17 270 20
rect 192 7 193 10
rect 195 7 203 10
rect 205 7 207 10
rect 219 9 225 15
rect 215 3 225 9
rect 260 15 270 17
rect 273 28 315 45
rect 273 27 293 28
rect 273 15 283 27
rect 288 26 291 27
rect 288 23 291 24
rect 299 24 315 28
rect 305 20 315 24
rect 301 17 302 20
rect 304 17 315 20
rect 237 7 238 10
rect 240 7 248 10
rect 250 7 252 10
rect 264 9 270 15
rect 260 3 270 9
rect 305 15 315 17
rect 318 28 360 45
rect 318 27 338 28
rect 318 15 328 27
rect 333 26 336 27
rect 333 23 336 24
rect 344 24 360 28
rect 350 20 360 24
rect 346 17 347 20
rect 349 17 360 20
rect 282 7 283 10
rect 285 7 293 10
rect 295 7 297 10
rect 309 9 315 15
rect 305 3 315 9
rect 350 15 360 17
rect 363 28 405 45
rect 363 27 383 28
rect 363 15 373 27
rect 378 26 381 27
rect 378 23 381 24
rect 389 24 405 28
rect 395 20 405 24
rect 391 17 392 20
rect 394 17 405 20
rect 327 7 328 10
rect 330 7 338 10
rect 340 7 342 10
rect 354 9 360 15
rect 350 3 360 9
rect 395 15 405 17
rect 408 28 450 45
rect 408 27 428 28
rect 408 15 418 27
rect 423 26 426 27
rect 423 23 426 24
rect 434 24 450 28
rect 440 20 450 24
rect 436 17 437 20
rect 439 17 450 20
rect 372 7 373 10
rect 375 7 383 10
rect 385 7 387 10
rect 399 9 405 15
rect 395 3 405 9
rect 440 15 450 17
rect 453 28 495 45
rect 453 27 473 28
rect 453 15 463 27
rect 468 26 471 27
rect 468 23 471 24
rect 479 24 495 28
rect 485 20 495 24
rect 481 17 482 20
rect 484 17 495 20
rect 417 7 418 10
rect 420 7 428 10
rect 430 7 432 10
rect 444 9 450 15
rect 440 3 450 9
rect 485 15 495 17
rect 498 28 540 45
rect 498 27 518 28
rect 498 15 508 27
rect 513 26 516 27
rect 513 23 516 24
rect 524 24 540 28
rect 530 20 540 24
rect 526 17 527 20
rect 529 17 540 20
rect 462 7 463 10
rect 465 7 473 10
rect 475 7 477 10
rect 489 9 495 15
rect 485 3 495 9
rect 530 15 540 17
rect 543 28 585 45
rect 543 27 563 28
rect 543 15 553 27
rect 558 26 561 27
rect 558 23 561 24
rect 569 24 585 28
rect 575 20 585 24
rect 571 17 572 20
rect 574 17 585 20
rect 507 7 508 10
rect 510 7 518 10
rect 520 7 522 10
rect 534 9 540 15
rect 530 3 540 9
rect 575 15 585 17
rect 588 28 630 45
rect 588 27 608 28
rect 588 15 598 27
rect 603 26 606 27
rect 603 23 606 24
rect 614 24 630 28
rect 620 20 630 24
rect 616 17 617 20
rect 619 17 630 20
rect 552 7 553 10
rect 555 7 563 10
rect 565 7 567 10
rect 579 9 585 15
rect 575 3 585 9
rect 620 15 630 17
rect 633 28 675 45
rect 633 27 653 28
rect 633 15 643 27
rect 648 26 651 27
rect 648 23 651 24
rect 659 24 675 28
rect 665 20 675 24
rect 661 17 662 20
rect 664 17 675 20
rect 597 7 598 10
rect 600 7 608 10
rect 610 7 612 10
rect 624 9 630 15
rect 620 3 630 9
rect 665 15 675 17
rect 678 28 720 45
rect 678 27 698 28
rect 678 15 688 27
rect 693 26 696 27
rect 693 23 696 24
rect 704 24 720 28
rect 710 20 720 24
rect 706 17 707 20
rect 709 17 720 20
rect 642 7 643 10
rect 645 7 653 10
rect 655 7 657 10
rect 669 9 675 15
rect 665 3 675 9
rect 710 15 720 17
rect 723 28 765 45
rect 723 27 743 28
rect 723 15 733 27
rect 738 26 741 27
rect 738 23 741 24
rect 749 24 765 28
rect 755 20 765 24
rect 751 17 752 20
rect 754 17 765 20
rect 687 7 688 10
rect 690 7 698 10
rect 700 7 702 10
rect 714 9 720 15
rect 710 3 720 9
rect 755 15 765 17
rect 768 28 810 45
rect 768 27 788 28
rect 768 15 778 27
rect 783 26 786 27
rect 783 23 786 24
rect 794 24 810 28
rect 800 20 810 24
rect 796 17 797 20
rect 799 17 810 20
rect 732 7 733 10
rect 735 7 743 10
rect 745 7 747 10
rect 759 9 765 15
rect 755 3 765 9
rect 800 15 810 17
rect 813 28 855 45
rect 813 27 833 28
rect 813 15 823 27
rect 828 26 831 27
rect 828 23 831 24
rect 839 24 855 28
rect 845 20 855 24
rect 841 17 842 20
rect 844 17 855 20
rect 777 7 778 10
rect 780 7 788 10
rect 790 7 792 10
rect 804 9 810 15
rect 800 3 810 9
rect 845 15 855 17
rect 858 28 900 45
rect 858 27 878 28
rect 858 15 868 27
rect 873 26 876 27
rect 873 23 876 24
rect 884 24 900 28
rect 890 20 900 24
rect 886 17 887 20
rect 889 17 900 20
rect 822 7 823 10
rect 825 7 833 10
rect 835 7 837 10
rect 849 9 855 15
rect 845 3 855 9
rect 890 15 900 17
rect 867 7 868 10
rect 870 7 878 10
rect 880 7 882 10
rect 894 9 900 15
rect 890 3 900 9
rect -213 -153 -171 -136
rect -213 -154 -193 -153
rect -268 -158 -263 -157
rect -268 -162 -266 -158
rect -268 -163 -263 -162
rect -298 -164 -292 -163
rect -298 -168 -297 -164
rect -293 -168 -292 -164
rect -298 -169 -292 -168
rect -290 -169 -287 -163
rect -285 -164 -280 -163
rect -285 -168 -284 -164
rect -285 -169 -280 -168
rect -268 -170 -263 -165
rect -213 -166 -203 -154
rect -198 -155 -195 -154
rect -198 -158 -195 -157
rect -187 -157 -171 -153
rect -181 -161 -171 -157
rect -185 -164 -184 -161
rect -182 -164 -171 -161
rect -268 -176 -260 -170
rect -258 -171 -253 -170
rect -258 -175 -257 -171
rect -181 -166 -171 -164
rect -204 -174 -203 -171
rect -201 -174 -193 -171
rect -191 -174 -189 -171
rect -177 -172 -171 -166
rect -258 -176 -253 -175
rect -268 -182 -262 -176
rect -181 -178 -171 -172
<< ndcontact >>
rect 17 874 21 878
rect 27 871 31 875
rect 8 862 12 866
rect 62 874 66 878
rect 72 871 76 875
rect 27 862 31 866
rect 53 862 57 866
rect 107 874 111 878
rect 117 871 121 875
rect 72 862 76 866
rect 98 862 102 866
rect 152 874 156 878
rect 162 871 166 875
rect 117 862 121 866
rect 143 862 147 866
rect 197 874 201 878
rect 207 871 211 875
rect 162 862 166 866
rect 188 862 192 866
rect 242 874 246 878
rect 252 871 256 875
rect 207 862 211 866
rect 233 862 237 866
rect 287 874 291 878
rect 297 871 301 875
rect 252 862 256 866
rect 278 862 282 866
rect 332 874 336 878
rect 342 871 346 875
rect 297 862 301 866
rect 323 862 327 866
rect 377 874 381 878
rect 387 871 391 875
rect 342 862 346 866
rect 368 862 372 866
rect 422 874 426 878
rect 432 871 436 875
rect 387 862 391 866
rect 413 862 417 866
rect 467 874 471 878
rect 477 871 481 875
rect 432 862 436 866
rect 458 862 462 866
rect 512 874 516 878
rect 522 871 526 875
rect 477 862 481 866
rect 503 862 507 866
rect 557 874 561 878
rect 567 871 571 875
rect 522 862 526 866
rect 548 862 552 866
rect 602 874 606 878
rect 612 871 616 875
rect 567 862 571 866
rect 593 862 597 866
rect 647 874 651 878
rect 657 871 661 875
rect 612 862 616 866
rect 638 862 642 866
rect 692 874 696 878
rect 702 871 706 875
rect 657 862 661 866
rect 683 862 687 866
rect 737 874 741 878
rect 747 871 751 875
rect 702 862 706 866
rect 728 862 732 866
rect 782 874 786 878
rect 792 871 796 875
rect 747 862 751 866
rect 773 862 777 866
rect 827 874 831 878
rect 837 871 841 875
rect 792 862 796 866
rect 818 862 822 866
rect 872 874 876 878
rect 882 871 886 875
rect 837 862 841 866
rect 863 862 867 866
rect 882 862 886 866
rect 17 829 21 833
rect 27 826 31 830
rect 8 817 12 821
rect 62 829 66 833
rect 72 826 76 830
rect 27 817 31 821
rect 53 817 57 821
rect 107 829 111 833
rect 117 826 121 830
rect 72 817 76 821
rect 98 817 102 821
rect 152 829 156 833
rect 162 826 166 830
rect 117 817 121 821
rect 143 817 147 821
rect 197 829 201 833
rect 207 826 211 830
rect 162 817 166 821
rect 188 817 192 821
rect 242 829 246 833
rect 252 826 256 830
rect 207 817 211 821
rect 233 817 237 821
rect 287 829 291 833
rect 297 826 301 830
rect 252 817 256 821
rect 278 817 282 821
rect 332 829 336 833
rect 342 826 346 830
rect 297 817 301 821
rect 323 817 327 821
rect 377 829 381 833
rect 387 826 391 830
rect 342 817 346 821
rect 368 817 372 821
rect 422 829 426 833
rect 432 826 436 830
rect 387 817 391 821
rect 413 817 417 821
rect 467 829 471 833
rect 477 826 481 830
rect 432 817 436 821
rect 458 817 462 821
rect 512 829 516 833
rect 522 826 526 830
rect 477 817 481 821
rect 503 817 507 821
rect 557 829 561 833
rect 567 826 571 830
rect 522 817 526 821
rect 548 817 552 821
rect 602 829 606 833
rect 612 826 616 830
rect 567 817 571 821
rect 593 817 597 821
rect 647 829 651 833
rect 657 826 661 830
rect 612 817 616 821
rect 638 817 642 821
rect 692 829 696 833
rect 702 826 706 830
rect 657 817 661 821
rect 683 817 687 821
rect 737 829 741 833
rect 747 826 751 830
rect 702 817 706 821
rect 728 817 732 821
rect 782 829 786 833
rect 792 826 796 830
rect 747 817 751 821
rect 773 817 777 821
rect 827 829 831 833
rect 837 826 841 830
rect 792 817 796 821
rect 818 817 822 821
rect 872 829 876 833
rect 882 826 886 830
rect 837 817 841 821
rect 863 817 867 821
rect 882 817 886 821
rect 17 784 21 788
rect 27 781 31 785
rect 8 772 12 776
rect 62 784 66 788
rect 72 781 76 785
rect 27 772 31 776
rect 53 772 57 776
rect 107 784 111 788
rect 117 781 121 785
rect 72 772 76 776
rect 98 772 102 776
rect 152 784 156 788
rect 162 781 166 785
rect 117 772 121 776
rect 143 772 147 776
rect 197 784 201 788
rect 207 781 211 785
rect 162 772 166 776
rect 188 772 192 776
rect 242 784 246 788
rect 252 781 256 785
rect 207 772 211 776
rect 233 772 237 776
rect 287 784 291 788
rect 297 781 301 785
rect 252 772 256 776
rect 278 772 282 776
rect 332 784 336 788
rect 342 781 346 785
rect 297 772 301 776
rect 323 772 327 776
rect 377 784 381 788
rect 387 781 391 785
rect 342 772 346 776
rect 368 772 372 776
rect 422 784 426 788
rect 432 781 436 785
rect 387 772 391 776
rect 413 772 417 776
rect 467 784 471 788
rect 477 781 481 785
rect 432 772 436 776
rect 458 772 462 776
rect 512 784 516 788
rect 522 781 526 785
rect 477 772 481 776
rect 503 772 507 776
rect 557 784 561 788
rect 567 781 571 785
rect 522 772 526 776
rect 548 772 552 776
rect 602 784 606 788
rect 612 781 616 785
rect 567 772 571 776
rect 593 772 597 776
rect 647 784 651 788
rect 657 781 661 785
rect 612 772 616 776
rect 638 772 642 776
rect 692 784 696 788
rect 702 781 706 785
rect 657 772 661 776
rect 683 772 687 776
rect 737 784 741 788
rect 747 781 751 785
rect 702 772 706 776
rect 728 772 732 776
rect 782 784 786 788
rect 792 781 796 785
rect 747 772 751 776
rect 773 772 777 776
rect 827 784 831 788
rect 837 781 841 785
rect 792 772 796 776
rect 818 772 822 776
rect 872 784 876 788
rect 882 781 886 785
rect 837 772 841 776
rect 863 772 867 776
rect 882 772 886 776
rect 17 739 21 743
rect 27 736 31 740
rect 8 727 12 731
rect 62 739 66 743
rect 72 736 76 740
rect 27 727 31 731
rect 53 727 57 731
rect 107 739 111 743
rect 117 736 121 740
rect 72 727 76 731
rect 98 727 102 731
rect 152 739 156 743
rect 162 736 166 740
rect 117 727 121 731
rect 143 727 147 731
rect 197 739 201 743
rect 207 736 211 740
rect 162 727 166 731
rect 188 727 192 731
rect 242 739 246 743
rect 252 736 256 740
rect 207 727 211 731
rect 233 727 237 731
rect 287 739 291 743
rect 297 736 301 740
rect 252 727 256 731
rect 278 727 282 731
rect 332 739 336 743
rect 342 736 346 740
rect 297 727 301 731
rect 323 727 327 731
rect 377 739 381 743
rect 387 736 391 740
rect 342 727 346 731
rect 368 727 372 731
rect 422 739 426 743
rect 432 736 436 740
rect 387 727 391 731
rect 413 727 417 731
rect 467 739 471 743
rect 477 736 481 740
rect 432 727 436 731
rect 458 727 462 731
rect 512 739 516 743
rect 522 736 526 740
rect 477 727 481 731
rect 503 727 507 731
rect 557 739 561 743
rect 567 736 571 740
rect 522 727 526 731
rect 548 727 552 731
rect 602 739 606 743
rect 612 736 616 740
rect 567 727 571 731
rect 593 727 597 731
rect 647 739 651 743
rect 657 736 661 740
rect 612 727 616 731
rect 638 727 642 731
rect 692 739 696 743
rect 702 736 706 740
rect 657 727 661 731
rect 683 727 687 731
rect 737 739 741 743
rect 747 736 751 740
rect 702 727 706 731
rect 728 727 732 731
rect 782 739 786 743
rect 792 736 796 740
rect 747 727 751 731
rect 773 727 777 731
rect 827 739 831 743
rect 837 736 841 740
rect 792 727 796 731
rect 818 727 822 731
rect 872 739 876 743
rect 882 736 886 740
rect 837 727 841 731
rect 863 727 867 731
rect 882 727 886 731
rect 17 694 21 698
rect 27 691 31 695
rect 8 682 12 686
rect 62 694 66 698
rect 72 691 76 695
rect 27 682 31 686
rect 53 682 57 686
rect 107 694 111 698
rect 117 691 121 695
rect 72 682 76 686
rect 98 682 102 686
rect 152 694 156 698
rect 162 691 166 695
rect 117 682 121 686
rect 143 682 147 686
rect 197 694 201 698
rect 207 691 211 695
rect 162 682 166 686
rect 188 682 192 686
rect 242 694 246 698
rect 252 691 256 695
rect 207 682 211 686
rect 233 682 237 686
rect 287 694 291 698
rect 297 691 301 695
rect 252 682 256 686
rect 278 682 282 686
rect 332 694 336 698
rect 342 691 346 695
rect 297 682 301 686
rect 323 682 327 686
rect 377 694 381 698
rect 387 691 391 695
rect 342 682 346 686
rect 368 682 372 686
rect 422 694 426 698
rect 432 691 436 695
rect 387 682 391 686
rect 413 682 417 686
rect 467 694 471 698
rect 477 691 481 695
rect 432 682 436 686
rect 458 682 462 686
rect 512 694 516 698
rect 522 691 526 695
rect 477 682 481 686
rect 503 682 507 686
rect 557 694 561 698
rect 567 691 571 695
rect 522 682 526 686
rect 548 682 552 686
rect 602 694 606 698
rect 612 691 616 695
rect 567 682 571 686
rect 593 682 597 686
rect 647 694 651 698
rect 657 691 661 695
rect 612 682 616 686
rect 638 682 642 686
rect 692 694 696 698
rect 702 691 706 695
rect 657 682 661 686
rect 683 682 687 686
rect 737 694 741 698
rect 747 691 751 695
rect 702 682 706 686
rect 728 682 732 686
rect 782 694 786 698
rect 792 691 796 695
rect 747 682 751 686
rect 773 682 777 686
rect 827 694 831 698
rect 837 691 841 695
rect 792 682 796 686
rect 818 682 822 686
rect 872 694 876 698
rect 882 691 886 695
rect 837 682 841 686
rect 863 682 867 686
rect 882 682 886 686
rect 17 649 21 653
rect 27 646 31 650
rect 8 637 12 641
rect 62 649 66 653
rect 72 646 76 650
rect 27 637 31 641
rect 53 637 57 641
rect 107 649 111 653
rect 117 646 121 650
rect 72 637 76 641
rect 98 637 102 641
rect 152 649 156 653
rect 162 646 166 650
rect 117 637 121 641
rect 143 637 147 641
rect 197 649 201 653
rect 207 646 211 650
rect 162 637 166 641
rect 188 637 192 641
rect 242 649 246 653
rect 252 646 256 650
rect 207 637 211 641
rect 233 637 237 641
rect 287 649 291 653
rect 297 646 301 650
rect 252 637 256 641
rect 278 637 282 641
rect 332 649 336 653
rect 342 646 346 650
rect 297 637 301 641
rect 323 637 327 641
rect 377 649 381 653
rect 387 646 391 650
rect 342 637 346 641
rect 368 637 372 641
rect 422 649 426 653
rect 432 646 436 650
rect 387 637 391 641
rect 413 637 417 641
rect 467 649 471 653
rect 477 646 481 650
rect 432 637 436 641
rect 458 637 462 641
rect 512 649 516 653
rect 522 646 526 650
rect 477 637 481 641
rect 503 637 507 641
rect 557 649 561 653
rect 567 646 571 650
rect 522 637 526 641
rect 548 637 552 641
rect 602 649 606 653
rect 612 646 616 650
rect 567 637 571 641
rect 593 637 597 641
rect 647 649 651 653
rect 657 646 661 650
rect 612 637 616 641
rect 638 637 642 641
rect 692 649 696 653
rect 702 646 706 650
rect 657 637 661 641
rect 683 637 687 641
rect 737 649 741 653
rect 747 646 751 650
rect 702 637 706 641
rect 728 637 732 641
rect 782 649 786 653
rect 792 646 796 650
rect 747 637 751 641
rect 773 637 777 641
rect 827 649 831 653
rect 837 646 841 650
rect 792 637 796 641
rect 818 637 822 641
rect 872 649 876 653
rect 882 646 886 650
rect 837 637 841 641
rect 863 637 867 641
rect 882 637 886 641
rect 17 604 21 608
rect 27 601 31 605
rect 8 592 12 596
rect 62 604 66 608
rect 72 601 76 605
rect 27 592 31 596
rect 53 592 57 596
rect 107 604 111 608
rect 117 601 121 605
rect 72 592 76 596
rect 98 592 102 596
rect 152 604 156 608
rect 162 601 166 605
rect 117 592 121 596
rect 143 592 147 596
rect 197 604 201 608
rect 207 601 211 605
rect 162 592 166 596
rect 188 592 192 596
rect 242 604 246 608
rect 252 601 256 605
rect 207 592 211 596
rect 233 592 237 596
rect 287 604 291 608
rect 297 601 301 605
rect 252 592 256 596
rect 278 592 282 596
rect 332 604 336 608
rect 342 601 346 605
rect 297 592 301 596
rect 323 592 327 596
rect 377 604 381 608
rect 387 601 391 605
rect 342 592 346 596
rect 368 592 372 596
rect 422 604 426 608
rect 432 601 436 605
rect 387 592 391 596
rect 413 592 417 596
rect 467 604 471 608
rect 477 601 481 605
rect 432 592 436 596
rect 458 592 462 596
rect 512 604 516 608
rect 522 601 526 605
rect 477 592 481 596
rect 503 592 507 596
rect 557 604 561 608
rect 567 601 571 605
rect 522 592 526 596
rect 548 592 552 596
rect 602 604 606 608
rect 612 601 616 605
rect 567 592 571 596
rect 593 592 597 596
rect 647 604 651 608
rect 657 601 661 605
rect 612 592 616 596
rect 638 592 642 596
rect 692 604 696 608
rect 702 601 706 605
rect 657 592 661 596
rect 683 592 687 596
rect 737 604 741 608
rect 747 601 751 605
rect 702 592 706 596
rect 728 592 732 596
rect 782 604 786 608
rect 792 601 796 605
rect 747 592 751 596
rect 773 592 777 596
rect 827 604 831 608
rect 837 601 841 605
rect 792 592 796 596
rect 818 592 822 596
rect 872 604 876 608
rect 882 601 886 605
rect 837 592 841 596
rect 863 592 867 596
rect 882 592 886 596
rect 17 559 21 563
rect 27 556 31 560
rect 8 547 12 551
rect 62 559 66 563
rect 72 556 76 560
rect 27 547 31 551
rect 53 547 57 551
rect 107 559 111 563
rect 117 556 121 560
rect 72 547 76 551
rect 98 547 102 551
rect 152 559 156 563
rect 162 556 166 560
rect 117 547 121 551
rect 143 547 147 551
rect 197 559 201 563
rect 207 556 211 560
rect 162 547 166 551
rect 188 547 192 551
rect 242 559 246 563
rect 252 556 256 560
rect 207 547 211 551
rect 233 547 237 551
rect 287 559 291 563
rect 297 556 301 560
rect 252 547 256 551
rect 278 547 282 551
rect 332 559 336 563
rect 342 556 346 560
rect 297 547 301 551
rect 323 547 327 551
rect 377 559 381 563
rect 387 556 391 560
rect 342 547 346 551
rect 368 547 372 551
rect 422 559 426 563
rect 432 556 436 560
rect 387 547 391 551
rect 413 547 417 551
rect 467 559 471 563
rect 477 556 481 560
rect 432 547 436 551
rect 458 547 462 551
rect 512 559 516 563
rect 522 556 526 560
rect 477 547 481 551
rect 503 547 507 551
rect 557 559 561 563
rect 567 556 571 560
rect 522 547 526 551
rect 548 547 552 551
rect 602 559 606 563
rect 612 556 616 560
rect 567 547 571 551
rect 593 547 597 551
rect 647 559 651 563
rect 657 556 661 560
rect 612 547 616 551
rect 638 547 642 551
rect 692 559 696 563
rect 702 556 706 560
rect 657 547 661 551
rect 683 547 687 551
rect 737 559 741 563
rect 747 556 751 560
rect 702 547 706 551
rect 728 547 732 551
rect 782 559 786 563
rect 792 556 796 560
rect 747 547 751 551
rect 773 547 777 551
rect 827 559 831 563
rect 837 556 841 560
rect 792 547 796 551
rect 818 547 822 551
rect 872 559 876 563
rect 882 556 886 560
rect 837 547 841 551
rect 863 547 867 551
rect 882 547 886 551
rect 17 514 21 518
rect 27 511 31 515
rect 8 502 12 506
rect 62 514 66 518
rect 72 511 76 515
rect 27 502 31 506
rect 53 502 57 506
rect 107 514 111 518
rect 117 511 121 515
rect 72 502 76 506
rect 98 502 102 506
rect 152 514 156 518
rect 162 511 166 515
rect 117 502 121 506
rect 143 502 147 506
rect 197 514 201 518
rect 207 511 211 515
rect 162 502 166 506
rect 188 502 192 506
rect 242 514 246 518
rect 252 511 256 515
rect 207 502 211 506
rect 233 502 237 506
rect 287 514 291 518
rect 297 511 301 515
rect 252 502 256 506
rect 278 502 282 506
rect 332 514 336 518
rect 342 511 346 515
rect 297 502 301 506
rect 323 502 327 506
rect 377 514 381 518
rect 387 511 391 515
rect 342 502 346 506
rect 368 502 372 506
rect 422 514 426 518
rect 432 511 436 515
rect 387 502 391 506
rect 413 502 417 506
rect 467 514 471 518
rect 477 511 481 515
rect 432 502 436 506
rect 458 502 462 506
rect 512 514 516 518
rect 522 511 526 515
rect 477 502 481 506
rect 503 502 507 506
rect 557 514 561 518
rect 567 511 571 515
rect 522 502 526 506
rect 548 502 552 506
rect 602 514 606 518
rect 612 511 616 515
rect 567 502 571 506
rect 593 502 597 506
rect 647 514 651 518
rect 657 511 661 515
rect 612 502 616 506
rect 638 502 642 506
rect 692 514 696 518
rect 702 511 706 515
rect 657 502 661 506
rect 683 502 687 506
rect 737 514 741 518
rect 747 511 751 515
rect 702 502 706 506
rect 728 502 732 506
rect 782 514 786 518
rect 792 511 796 515
rect 747 502 751 506
rect 773 502 777 506
rect 827 514 831 518
rect 837 511 841 515
rect 792 502 796 506
rect 818 502 822 506
rect 872 514 876 518
rect 882 511 886 515
rect 837 502 841 506
rect 863 502 867 506
rect 882 502 886 506
rect 17 469 21 473
rect 27 466 31 470
rect 8 457 12 461
rect 62 469 66 473
rect 72 466 76 470
rect 27 457 31 461
rect 53 457 57 461
rect 107 469 111 473
rect 117 466 121 470
rect 72 457 76 461
rect 98 457 102 461
rect 152 469 156 473
rect 162 466 166 470
rect 117 457 121 461
rect 143 457 147 461
rect 197 469 201 473
rect 207 466 211 470
rect 162 457 166 461
rect 188 457 192 461
rect 242 469 246 473
rect 252 466 256 470
rect 207 457 211 461
rect 233 457 237 461
rect 287 469 291 473
rect 297 466 301 470
rect 252 457 256 461
rect 278 457 282 461
rect 332 469 336 473
rect 342 466 346 470
rect 297 457 301 461
rect 323 457 327 461
rect 377 469 381 473
rect 387 466 391 470
rect 342 457 346 461
rect 368 457 372 461
rect 422 469 426 473
rect 432 466 436 470
rect 387 457 391 461
rect 413 457 417 461
rect 467 469 471 473
rect 477 466 481 470
rect 432 457 436 461
rect 458 457 462 461
rect 512 469 516 473
rect 522 466 526 470
rect 477 457 481 461
rect 503 457 507 461
rect 557 469 561 473
rect 567 466 571 470
rect 522 457 526 461
rect 548 457 552 461
rect 602 469 606 473
rect 612 466 616 470
rect 567 457 571 461
rect 593 457 597 461
rect 647 469 651 473
rect 657 466 661 470
rect 612 457 616 461
rect 638 457 642 461
rect 692 469 696 473
rect 702 466 706 470
rect 657 457 661 461
rect 683 457 687 461
rect 737 469 741 473
rect 747 466 751 470
rect 702 457 706 461
rect 728 457 732 461
rect 782 469 786 473
rect 792 466 796 470
rect 747 457 751 461
rect 773 457 777 461
rect 827 469 831 473
rect 837 466 841 470
rect 792 457 796 461
rect 818 457 822 461
rect 872 469 876 473
rect 882 466 886 470
rect 837 457 841 461
rect 863 457 867 461
rect 882 457 886 461
rect 17 424 21 428
rect 27 421 31 425
rect 8 412 12 416
rect 62 424 66 428
rect 72 421 76 425
rect 27 412 31 416
rect 53 412 57 416
rect 107 424 111 428
rect 117 421 121 425
rect 72 412 76 416
rect 98 412 102 416
rect 152 424 156 428
rect 162 421 166 425
rect 117 412 121 416
rect 143 412 147 416
rect 197 424 201 428
rect 207 421 211 425
rect 162 412 166 416
rect 188 412 192 416
rect 242 424 246 428
rect 252 421 256 425
rect 207 412 211 416
rect 233 412 237 416
rect 287 424 291 428
rect 297 421 301 425
rect 252 412 256 416
rect 278 412 282 416
rect 332 424 336 428
rect 342 421 346 425
rect 297 412 301 416
rect 323 412 327 416
rect 377 424 381 428
rect 387 421 391 425
rect 342 412 346 416
rect 368 412 372 416
rect 422 424 426 428
rect 432 421 436 425
rect 387 412 391 416
rect 413 412 417 416
rect 467 424 471 428
rect 477 421 481 425
rect 432 412 436 416
rect 458 412 462 416
rect 512 424 516 428
rect 522 421 526 425
rect 477 412 481 416
rect 503 412 507 416
rect 557 424 561 428
rect 567 421 571 425
rect 522 412 526 416
rect 548 412 552 416
rect 602 424 606 428
rect 612 421 616 425
rect 567 412 571 416
rect 593 412 597 416
rect 647 424 651 428
rect 657 421 661 425
rect 612 412 616 416
rect 638 412 642 416
rect 692 424 696 428
rect 702 421 706 425
rect 657 412 661 416
rect 683 412 687 416
rect 737 424 741 428
rect 747 421 751 425
rect 702 412 706 416
rect 728 412 732 416
rect 782 424 786 428
rect 792 421 796 425
rect 747 412 751 416
rect 773 412 777 416
rect 827 424 831 428
rect 837 421 841 425
rect 792 412 796 416
rect 818 412 822 416
rect 872 424 876 428
rect 882 421 886 425
rect 837 412 841 416
rect 863 412 867 416
rect 882 412 886 416
rect 17 379 21 383
rect 27 376 31 380
rect 8 367 12 371
rect 62 379 66 383
rect 72 376 76 380
rect 27 367 31 371
rect 53 367 57 371
rect 107 379 111 383
rect 117 376 121 380
rect 72 367 76 371
rect 98 367 102 371
rect 152 379 156 383
rect 162 376 166 380
rect 117 367 121 371
rect 143 367 147 371
rect 197 379 201 383
rect 207 376 211 380
rect 162 367 166 371
rect 188 367 192 371
rect 242 379 246 383
rect 252 376 256 380
rect 207 367 211 371
rect 233 367 237 371
rect 287 379 291 383
rect 297 376 301 380
rect 252 367 256 371
rect 278 367 282 371
rect 332 379 336 383
rect 342 376 346 380
rect 297 367 301 371
rect 323 367 327 371
rect 377 379 381 383
rect 387 376 391 380
rect 342 367 346 371
rect 368 367 372 371
rect 422 379 426 383
rect 432 376 436 380
rect 387 367 391 371
rect 413 367 417 371
rect 467 379 471 383
rect 477 376 481 380
rect 432 367 436 371
rect 458 367 462 371
rect 512 379 516 383
rect 522 376 526 380
rect 477 367 481 371
rect 503 367 507 371
rect 557 379 561 383
rect 567 376 571 380
rect 522 367 526 371
rect 548 367 552 371
rect 602 379 606 383
rect 612 376 616 380
rect 567 367 571 371
rect 593 367 597 371
rect 647 379 651 383
rect 657 376 661 380
rect 612 367 616 371
rect 638 367 642 371
rect 692 379 696 383
rect 702 376 706 380
rect 657 367 661 371
rect 683 367 687 371
rect 737 379 741 383
rect 747 376 751 380
rect 702 367 706 371
rect 728 367 732 371
rect 782 379 786 383
rect 792 376 796 380
rect 747 367 751 371
rect 773 367 777 371
rect 827 379 831 383
rect 837 376 841 380
rect 792 367 796 371
rect 818 367 822 371
rect 872 379 876 383
rect 882 376 886 380
rect 837 367 841 371
rect 863 367 867 371
rect 882 367 886 371
rect 17 334 21 338
rect 27 331 31 335
rect 8 322 12 326
rect 62 334 66 338
rect 72 331 76 335
rect 27 322 31 326
rect 53 322 57 326
rect 107 334 111 338
rect 117 331 121 335
rect 72 322 76 326
rect 98 322 102 326
rect 152 334 156 338
rect 162 331 166 335
rect 117 322 121 326
rect 143 322 147 326
rect 197 334 201 338
rect 207 331 211 335
rect 162 322 166 326
rect 188 322 192 326
rect 242 334 246 338
rect 252 331 256 335
rect 207 322 211 326
rect 233 322 237 326
rect 287 334 291 338
rect 297 331 301 335
rect 252 322 256 326
rect 278 322 282 326
rect 332 334 336 338
rect 342 331 346 335
rect 297 322 301 326
rect 323 322 327 326
rect 377 334 381 338
rect 387 331 391 335
rect 342 322 346 326
rect 368 322 372 326
rect 422 334 426 338
rect 432 331 436 335
rect 387 322 391 326
rect 413 322 417 326
rect 467 334 471 338
rect 477 331 481 335
rect 432 322 436 326
rect 458 322 462 326
rect 512 334 516 338
rect 522 331 526 335
rect 477 322 481 326
rect 503 322 507 326
rect 557 334 561 338
rect 567 331 571 335
rect 522 322 526 326
rect 548 322 552 326
rect 602 334 606 338
rect 612 331 616 335
rect 567 322 571 326
rect 593 322 597 326
rect 647 334 651 338
rect 657 331 661 335
rect 612 322 616 326
rect 638 322 642 326
rect 692 334 696 338
rect 702 331 706 335
rect 657 322 661 326
rect 683 322 687 326
rect 737 334 741 338
rect 747 331 751 335
rect 702 322 706 326
rect 728 322 732 326
rect 782 334 786 338
rect 792 331 796 335
rect 747 322 751 326
rect 773 322 777 326
rect 827 334 831 338
rect 837 331 841 335
rect 792 322 796 326
rect 818 322 822 326
rect 872 334 876 338
rect 882 331 886 335
rect 837 322 841 326
rect 863 322 867 326
rect 882 322 886 326
rect 17 289 21 293
rect 27 286 31 290
rect 8 277 12 281
rect 62 289 66 293
rect 72 286 76 290
rect 27 277 31 281
rect 53 277 57 281
rect 107 289 111 293
rect 117 286 121 290
rect 72 277 76 281
rect 98 277 102 281
rect 152 289 156 293
rect 162 286 166 290
rect 117 277 121 281
rect 143 277 147 281
rect 197 289 201 293
rect 207 286 211 290
rect 162 277 166 281
rect 188 277 192 281
rect 242 289 246 293
rect 252 286 256 290
rect 207 277 211 281
rect 233 277 237 281
rect 287 289 291 293
rect 297 286 301 290
rect 252 277 256 281
rect 278 277 282 281
rect 332 289 336 293
rect 342 286 346 290
rect 297 277 301 281
rect 323 277 327 281
rect 377 289 381 293
rect 387 286 391 290
rect 342 277 346 281
rect 368 277 372 281
rect 422 289 426 293
rect 432 286 436 290
rect 387 277 391 281
rect 413 277 417 281
rect 467 289 471 293
rect 477 286 481 290
rect 432 277 436 281
rect 458 277 462 281
rect 512 289 516 293
rect 522 286 526 290
rect 477 277 481 281
rect 503 277 507 281
rect 557 289 561 293
rect 567 286 571 290
rect 522 277 526 281
rect 548 277 552 281
rect 602 289 606 293
rect 612 286 616 290
rect 567 277 571 281
rect 593 277 597 281
rect 647 289 651 293
rect 657 286 661 290
rect 612 277 616 281
rect 638 277 642 281
rect 692 289 696 293
rect 702 286 706 290
rect 657 277 661 281
rect 683 277 687 281
rect 737 289 741 293
rect 747 286 751 290
rect 702 277 706 281
rect 728 277 732 281
rect 782 289 786 293
rect 792 286 796 290
rect 747 277 751 281
rect 773 277 777 281
rect 827 289 831 293
rect 837 286 841 290
rect 792 277 796 281
rect 818 277 822 281
rect 872 289 876 293
rect 882 286 886 290
rect 837 277 841 281
rect 863 277 867 281
rect 882 277 886 281
rect 17 244 21 248
rect 27 241 31 245
rect 8 232 12 236
rect 62 244 66 248
rect 72 241 76 245
rect 27 232 31 236
rect 53 232 57 236
rect 107 244 111 248
rect 117 241 121 245
rect 72 232 76 236
rect 98 232 102 236
rect 152 244 156 248
rect 162 241 166 245
rect 117 232 121 236
rect 143 232 147 236
rect 197 244 201 248
rect 207 241 211 245
rect 162 232 166 236
rect 188 232 192 236
rect 242 244 246 248
rect 252 241 256 245
rect 207 232 211 236
rect 233 232 237 236
rect 287 244 291 248
rect 297 241 301 245
rect 252 232 256 236
rect 278 232 282 236
rect 332 244 336 248
rect 342 241 346 245
rect 297 232 301 236
rect 323 232 327 236
rect 377 244 381 248
rect 387 241 391 245
rect 342 232 346 236
rect 368 232 372 236
rect 422 244 426 248
rect 432 241 436 245
rect 387 232 391 236
rect 413 232 417 236
rect 467 244 471 248
rect 477 241 481 245
rect 432 232 436 236
rect 458 232 462 236
rect 512 244 516 248
rect 522 241 526 245
rect 477 232 481 236
rect 503 232 507 236
rect 557 244 561 248
rect 567 241 571 245
rect 522 232 526 236
rect 548 232 552 236
rect 602 244 606 248
rect 612 241 616 245
rect 567 232 571 236
rect 593 232 597 236
rect 647 244 651 248
rect 657 241 661 245
rect 612 232 616 236
rect 638 232 642 236
rect 692 244 696 248
rect 702 241 706 245
rect 657 232 661 236
rect 683 232 687 236
rect 737 244 741 248
rect 747 241 751 245
rect 702 232 706 236
rect 728 232 732 236
rect 782 244 786 248
rect 792 241 796 245
rect 747 232 751 236
rect 773 232 777 236
rect 827 244 831 248
rect 837 241 841 245
rect 792 232 796 236
rect 818 232 822 236
rect 872 244 876 248
rect 882 241 886 245
rect 837 232 841 236
rect 863 232 867 236
rect 882 232 886 236
rect 17 199 21 203
rect 27 196 31 200
rect 8 187 12 191
rect 62 199 66 203
rect 72 196 76 200
rect 27 187 31 191
rect 53 187 57 191
rect 107 199 111 203
rect 117 196 121 200
rect 72 187 76 191
rect 98 187 102 191
rect 152 199 156 203
rect 162 196 166 200
rect 117 187 121 191
rect 143 187 147 191
rect 197 199 201 203
rect 207 196 211 200
rect 162 187 166 191
rect 188 187 192 191
rect 242 199 246 203
rect 252 196 256 200
rect 207 187 211 191
rect 233 187 237 191
rect 287 199 291 203
rect 297 196 301 200
rect 252 187 256 191
rect 278 187 282 191
rect 332 199 336 203
rect 342 196 346 200
rect 297 187 301 191
rect 323 187 327 191
rect 377 199 381 203
rect 387 196 391 200
rect 342 187 346 191
rect 368 187 372 191
rect 422 199 426 203
rect 432 196 436 200
rect 387 187 391 191
rect 413 187 417 191
rect 467 199 471 203
rect 477 196 481 200
rect 432 187 436 191
rect 458 187 462 191
rect 512 199 516 203
rect 522 196 526 200
rect 477 187 481 191
rect 503 187 507 191
rect 557 199 561 203
rect 567 196 571 200
rect 522 187 526 191
rect 548 187 552 191
rect 602 199 606 203
rect 612 196 616 200
rect 567 187 571 191
rect 593 187 597 191
rect 647 199 651 203
rect 657 196 661 200
rect 612 187 616 191
rect 638 187 642 191
rect 692 199 696 203
rect 702 196 706 200
rect 657 187 661 191
rect 683 187 687 191
rect 737 199 741 203
rect 747 196 751 200
rect 702 187 706 191
rect 728 187 732 191
rect 782 199 786 203
rect 792 196 796 200
rect 747 187 751 191
rect 773 187 777 191
rect 827 199 831 203
rect 837 196 841 200
rect 792 187 796 191
rect 818 187 822 191
rect 872 199 876 203
rect 882 196 886 200
rect 837 187 841 191
rect 863 187 867 191
rect 882 187 886 191
rect 17 154 21 158
rect 27 151 31 155
rect 8 142 12 146
rect 62 154 66 158
rect 72 151 76 155
rect 27 142 31 146
rect 53 142 57 146
rect 107 154 111 158
rect 117 151 121 155
rect 72 142 76 146
rect 98 142 102 146
rect 152 154 156 158
rect 162 151 166 155
rect 117 142 121 146
rect 143 142 147 146
rect 197 154 201 158
rect 207 151 211 155
rect 162 142 166 146
rect 188 142 192 146
rect 242 154 246 158
rect 252 151 256 155
rect 207 142 211 146
rect 233 142 237 146
rect 287 154 291 158
rect 297 151 301 155
rect 252 142 256 146
rect 278 142 282 146
rect 332 154 336 158
rect 342 151 346 155
rect 297 142 301 146
rect 323 142 327 146
rect 377 154 381 158
rect 387 151 391 155
rect 342 142 346 146
rect 368 142 372 146
rect 422 154 426 158
rect 432 151 436 155
rect 387 142 391 146
rect 413 142 417 146
rect 467 154 471 158
rect 477 151 481 155
rect 432 142 436 146
rect 458 142 462 146
rect 512 154 516 158
rect 522 151 526 155
rect 477 142 481 146
rect 503 142 507 146
rect 557 154 561 158
rect 567 151 571 155
rect 522 142 526 146
rect 548 142 552 146
rect 602 154 606 158
rect 612 151 616 155
rect 567 142 571 146
rect 593 142 597 146
rect 647 154 651 158
rect 657 151 661 155
rect 612 142 616 146
rect 638 142 642 146
rect 692 154 696 158
rect 702 151 706 155
rect 657 142 661 146
rect 683 142 687 146
rect 737 154 741 158
rect 747 151 751 155
rect 702 142 706 146
rect 728 142 732 146
rect 782 154 786 158
rect 792 151 796 155
rect 747 142 751 146
rect 773 142 777 146
rect 827 154 831 158
rect 837 151 841 155
rect 792 142 796 146
rect 818 142 822 146
rect 872 154 876 158
rect 882 151 886 155
rect 837 142 841 146
rect 863 142 867 146
rect 882 142 886 146
rect 17 109 21 113
rect 27 106 31 110
rect 8 97 12 101
rect 62 109 66 113
rect 72 106 76 110
rect 27 97 31 101
rect 53 97 57 101
rect 107 109 111 113
rect 117 106 121 110
rect 72 97 76 101
rect 98 97 102 101
rect 152 109 156 113
rect 162 106 166 110
rect 117 97 121 101
rect 143 97 147 101
rect 197 109 201 113
rect 207 106 211 110
rect 162 97 166 101
rect 188 97 192 101
rect 242 109 246 113
rect 252 106 256 110
rect 207 97 211 101
rect 233 97 237 101
rect 287 109 291 113
rect 297 106 301 110
rect 252 97 256 101
rect 278 97 282 101
rect 332 109 336 113
rect 342 106 346 110
rect 297 97 301 101
rect 323 97 327 101
rect 377 109 381 113
rect 387 106 391 110
rect 342 97 346 101
rect 368 97 372 101
rect 422 109 426 113
rect 432 106 436 110
rect 387 97 391 101
rect 413 97 417 101
rect 467 109 471 113
rect 477 106 481 110
rect 432 97 436 101
rect 458 97 462 101
rect 512 109 516 113
rect 522 106 526 110
rect 477 97 481 101
rect 503 97 507 101
rect 557 109 561 113
rect 567 106 571 110
rect 522 97 526 101
rect 548 97 552 101
rect 602 109 606 113
rect 612 106 616 110
rect 567 97 571 101
rect 593 97 597 101
rect 647 109 651 113
rect 657 106 661 110
rect 612 97 616 101
rect 638 97 642 101
rect 692 109 696 113
rect 702 106 706 110
rect 657 97 661 101
rect 683 97 687 101
rect 737 109 741 113
rect 747 106 751 110
rect 702 97 706 101
rect 728 97 732 101
rect 782 109 786 113
rect 792 106 796 110
rect 747 97 751 101
rect 773 97 777 101
rect 827 109 831 113
rect 837 106 841 110
rect 792 97 796 101
rect 818 97 822 101
rect 872 109 876 113
rect 882 106 886 110
rect 837 97 841 101
rect 863 97 867 101
rect 882 97 886 101
rect 17 64 21 68
rect 27 61 31 65
rect 8 52 12 56
rect 62 64 66 68
rect 72 61 76 65
rect 27 52 31 56
rect 53 52 57 56
rect 107 64 111 68
rect 117 61 121 65
rect 72 52 76 56
rect 98 52 102 56
rect 152 64 156 68
rect 162 61 166 65
rect 117 52 121 56
rect 143 52 147 56
rect 197 64 201 68
rect 207 61 211 65
rect 162 52 166 56
rect 188 52 192 56
rect 242 64 246 68
rect 252 61 256 65
rect 207 52 211 56
rect 233 52 237 56
rect 287 64 291 68
rect 297 61 301 65
rect 252 52 256 56
rect 278 52 282 56
rect 332 64 336 68
rect 342 61 346 65
rect 297 52 301 56
rect 323 52 327 56
rect 377 64 381 68
rect 387 61 391 65
rect 342 52 346 56
rect 368 52 372 56
rect 422 64 426 68
rect 432 61 436 65
rect 387 52 391 56
rect 413 52 417 56
rect 467 64 471 68
rect 477 61 481 65
rect 432 52 436 56
rect 458 52 462 56
rect 512 64 516 68
rect 522 61 526 65
rect 477 52 481 56
rect 503 52 507 56
rect 557 64 561 68
rect 567 61 571 65
rect 522 52 526 56
rect 548 52 552 56
rect 602 64 606 68
rect 612 61 616 65
rect 567 52 571 56
rect 593 52 597 56
rect 647 64 651 68
rect 657 61 661 65
rect 612 52 616 56
rect 638 52 642 56
rect 692 64 696 68
rect 702 61 706 65
rect 657 52 661 56
rect 683 52 687 56
rect 737 64 741 68
rect 747 61 751 65
rect 702 52 706 56
rect 728 52 732 56
rect 782 64 786 68
rect 792 61 796 65
rect 747 52 751 56
rect 773 52 777 56
rect 827 64 831 68
rect 837 61 841 65
rect 792 52 796 56
rect 818 52 822 56
rect 872 64 876 68
rect 882 61 886 65
rect 837 52 841 56
rect 863 52 867 56
rect 882 52 886 56
rect 17 19 21 23
rect 27 16 31 20
rect 8 7 12 11
rect 62 19 66 23
rect 72 16 76 20
rect 27 7 31 11
rect 53 7 57 11
rect 107 19 111 23
rect 117 16 121 20
rect 72 7 76 11
rect 98 7 102 11
rect 152 19 156 23
rect 162 16 166 20
rect 117 7 121 11
rect 143 7 147 11
rect 197 19 201 23
rect 207 16 211 20
rect 162 7 166 11
rect 188 7 192 11
rect 242 19 246 23
rect 252 16 256 20
rect 207 7 211 11
rect 233 7 237 11
rect 287 19 291 23
rect 297 16 301 20
rect 252 7 256 11
rect 278 7 282 11
rect 332 19 336 23
rect 342 16 346 20
rect 297 7 301 11
rect 323 7 327 11
rect 377 19 381 23
rect 387 16 391 20
rect 342 7 346 11
rect 368 7 372 11
rect 422 19 426 23
rect 432 16 436 20
rect 387 7 391 11
rect 413 7 417 11
rect 467 19 471 23
rect 477 16 481 20
rect 432 7 436 11
rect 458 7 462 11
rect 512 19 516 23
rect 522 16 526 20
rect 477 7 481 11
rect 503 7 507 11
rect 557 19 561 23
rect 567 16 571 20
rect 522 7 526 11
rect 548 7 552 11
rect 602 19 606 23
rect 612 16 616 20
rect 567 7 571 11
rect 593 7 597 11
rect 647 19 651 23
rect 657 16 661 20
rect 612 7 616 11
rect 638 7 642 11
rect 692 19 696 23
rect 702 16 706 20
rect 657 7 661 11
rect 683 7 687 11
rect 737 19 741 23
rect 747 16 751 20
rect 702 7 706 11
rect 728 7 732 11
rect 782 19 786 23
rect 792 16 796 20
rect 747 7 751 11
rect 773 7 777 11
rect 827 19 831 23
rect 837 16 841 20
rect 792 7 796 11
rect 818 7 822 11
rect 872 19 876 23
rect 882 16 886 20
rect 837 7 841 11
rect 863 7 867 11
rect 882 7 886 11
rect -266 -162 -262 -158
rect -297 -168 -293 -164
rect -284 -168 -280 -164
rect -199 -162 -195 -158
rect -189 -165 -185 -161
rect -257 -175 -253 -171
rect -208 -174 -204 -170
rect -189 -174 -185 -170
<< polysilicon >>
rect 16 879 18 881
rect 21 879 24 881
rect 32 875 34 877
rect 13 865 15 867
rect 23 865 25 869
rect 32 866 34 872
rect 61 879 63 881
rect 66 879 69 881
rect 77 875 79 877
rect 13 857 15 862
rect 23 860 25 862
rect 58 865 60 867
rect 68 865 70 869
rect 77 866 79 872
rect 106 879 108 881
rect 111 879 114 881
rect 122 875 124 877
rect 58 857 60 862
rect 68 860 70 862
rect 103 865 105 867
rect 113 865 115 869
rect 122 866 124 872
rect 151 879 153 881
rect 156 879 159 881
rect 167 875 169 877
rect 103 857 105 862
rect 113 860 115 862
rect 148 865 150 867
rect 158 865 160 869
rect 167 866 169 872
rect 196 879 198 881
rect 201 879 204 881
rect 212 875 214 877
rect 148 857 150 862
rect 158 860 160 862
rect 193 865 195 867
rect 203 865 205 869
rect 212 866 214 872
rect 241 879 243 881
rect 246 879 249 881
rect 257 875 259 877
rect 193 857 195 862
rect 203 860 205 862
rect 238 865 240 867
rect 248 865 250 869
rect 257 866 259 872
rect 286 879 288 881
rect 291 879 294 881
rect 302 875 304 877
rect 238 857 240 862
rect 248 860 250 862
rect 283 865 285 867
rect 293 865 295 869
rect 302 866 304 872
rect 331 879 333 881
rect 336 879 339 881
rect 347 875 349 877
rect 283 857 285 862
rect 293 860 295 862
rect 328 865 330 867
rect 338 865 340 869
rect 347 866 349 872
rect 376 879 378 881
rect 381 879 384 881
rect 392 875 394 877
rect 328 857 330 862
rect 338 860 340 862
rect 373 865 375 867
rect 383 865 385 869
rect 392 866 394 872
rect 421 879 423 881
rect 426 879 429 881
rect 437 875 439 877
rect 373 857 375 862
rect 383 860 385 862
rect 418 865 420 867
rect 428 865 430 869
rect 437 866 439 872
rect 466 879 468 881
rect 471 879 474 881
rect 482 875 484 877
rect 418 857 420 862
rect 428 860 430 862
rect 463 865 465 867
rect 473 865 475 869
rect 482 866 484 872
rect 511 879 513 881
rect 516 879 519 881
rect 527 875 529 877
rect 463 857 465 862
rect 473 860 475 862
rect 508 865 510 867
rect 518 865 520 869
rect 527 866 529 872
rect 556 879 558 881
rect 561 879 564 881
rect 572 875 574 877
rect 508 857 510 862
rect 518 860 520 862
rect 553 865 555 867
rect 563 865 565 869
rect 572 866 574 872
rect 601 879 603 881
rect 606 879 609 881
rect 617 875 619 877
rect 553 857 555 862
rect 563 860 565 862
rect 598 865 600 867
rect 608 865 610 869
rect 617 866 619 872
rect 646 879 648 881
rect 651 879 654 881
rect 662 875 664 877
rect 598 857 600 862
rect 608 860 610 862
rect 643 865 645 867
rect 653 865 655 869
rect 662 866 664 872
rect 691 879 693 881
rect 696 879 699 881
rect 707 875 709 877
rect 643 857 645 862
rect 653 860 655 862
rect 688 865 690 867
rect 698 865 700 869
rect 707 866 709 872
rect 736 879 738 881
rect 741 879 744 881
rect 752 875 754 877
rect 688 857 690 862
rect 698 860 700 862
rect 733 865 735 867
rect 743 865 745 869
rect 752 866 754 872
rect 781 879 783 881
rect 786 879 789 881
rect 797 875 799 877
rect 733 857 735 862
rect 743 860 745 862
rect 778 865 780 867
rect 788 865 790 869
rect 797 866 799 872
rect 826 879 828 881
rect 831 879 834 881
rect 842 875 844 877
rect 778 857 780 862
rect 788 860 790 862
rect 823 865 825 867
rect 833 865 835 869
rect 842 866 844 872
rect 871 879 873 881
rect 876 879 879 881
rect 887 875 889 877
rect 823 857 825 862
rect 833 860 835 862
rect 868 865 870 867
rect 878 865 880 869
rect 887 866 889 872
rect 868 857 870 862
rect 878 860 880 862
rect 16 834 18 836
rect 21 834 24 836
rect 32 830 34 832
rect 13 820 15 822
rect 23 820 25 824
rect 32 821 34 827
rect 61 834 63 836
rect 66 834 69 836
rect 77 830 79 832
rect 13 812 15 817
rect 23 815 25 817
rect 58 820 60 822
rect 68 820 70 824
rect 77 821 79 827
rect 106 834 108 836
rect 111 834 114 836
rect 122 830 124 832
rect 58 812 60 817
rect 68 815 70 817
rect 103 820 105 822
rect 113 820 115 824
rect 122 821 124 827
rect 151 834 153 836
rect 156 834 159 836
rect 167 830 169 832
rect 103 812 105 817
rect 113 815 115 817
rect 148 820 150 822
rect 158 820 160 824
rect 167 821 169 827
rect 196 834 198 836
rect 201 834 204 836
rect 212 830 214 832
rect 148 812 150 817
rect 158 815 160 817
rect 193 820 195 822
rect 203 820 205 824
rect 212 821 214 827
rect 241 834 243 836
rect 246 834 249 836
rect 257 830 259 832
rect 193 812 195 817
rect 203 815 205 817
rect 238 820 240 822
rect 248 820 250 824
rect 257 821 259 827
rect 286 834 288 836
rect 291 834 294 836
rect 302 830 304 832
rect 238 812 240 817
rect 248 815 250 817
rect 283 820 285 822
rect 293 820 295 824
rect 302 821 304 827
rect 331 834 333 836
rect 336 834 339 836
rect 347 830 349 832
rect 283 812 285 817
rect 293 815 295 817
rect 328 820 330 822
rect 338 820 340 824
rect 347 821 349 827
rect 376 834 378 836
rect 381 834 384 836
rect 392 830 394 832
rect 328 812 330 817
rect 338 815 340 817
rect 373 820 375 822
rect 383 820 385 824
rect 392 821 394 827
rect 421 834 423 836
rect 426 834 429 836
rect 437 830 439 832
rect 373 812 375 817
rect 383 815 385 817
rect 418 820 420 822
rect 428 820 430 824
rect 437 821 439 827
rect 466 834 468 836
rect 471 834 474 836
rect 482 830 484 832
rect 418 812 420 817
rect 428 815 430 817
rect 463 820 465 822
rect 473 820 475 824
rect 482 821 484 827
rect 511 834 513 836
rect 516 834 519 836
rect 527 830 529 832
rect 463 812 465 817
rect 473 815 475 817
rect 508 820 510 822
rect 518 820 520 824
rect 527 821 529 827
rect 556 834 558 836
rect 561 834 564 836
rect 572 830 574 832
rect 508 812 510 817
rect 518 815 520 817
rect 553 820 555 822
rect 563 820 565 824
rect 572 821 574 827
rect 601 834 603 836
rect 606 834 609 836
rect 617 830 619 832
rect 553 812 555 817
rect 563 815 565 817
rect 598 820 600 822
rect 608 820 610 824
rect 617 821 619 827
rect 646 834 648 836
rect 651 834 654 836
rect 662 830 664 832
rect 598 812 600 817
rect 608 815 610 817
rect 643 820 645 822
rect 653 820 655 824
rect 662 821 664 827
rect 691 834 693 836
rect 696 834 699 836
rect 707 830 709 832
rect 643 812 645 817
rect 653 815 655 817
rect 688 820 690 822
rect 698 820 700 824
rect 707 821 709 827
rect 736 834 738 836
rect 741 834 744 836
rect 752 830 754 832
rect 688 812 690 817
rect 698 815 700 817
rect 733 820 735 822
rect 743 820 745 824
rect 752 821 754 827
rect 781 834 783 836
rect 786 834 789 836
rect 797 830 799 832
rect 733 812 735 817
rect 743 815 745 817
rect 778 820 780 822
rect 788 820 790 824
rect 797 821 799 827
rect 826 834 828 836
rect 831 834 834 836
rect 842 830 844 832
rect 778 812 780 817
rect 788 815 790 817
rect 823 820 825 822
rect 833 820 835 824
rect 842 821 844 827
rect 871 834 873 836
rect 876 834 879 836
rect 887 830 889 832
rect 823 812 825 817
rect 833 815 835 817
rect 868 820 870 822
rect 878 820 880 824
rect 887 821 889 827
rect 868 812 870 817
rect 878 815 880 817
rect 16 789 18 791
rect 21 789 24 791
rect 32 785 34 787
rect 13 775 15 777
rect 23 775 25 779
rect 32 776 34 782
rect 61 789 63 791
rect 66 789 69 791
rect 77 785 79 787
rect 13 767 15 772
rect 23 770 25 772
rect 58 775 60 777
rect 68 775 70 779
rect 77 776 79 782
rect 106 789 108 791
rect 111 789 114 791
rect 122 785 124 787
rect 58 767 60 772
rect 68 770 70 772
rect 103 775 105 777
rect 113 775 115 779
rect 122 776 124 782
rect 151 789 153 791
rect 156 789 159 791
rect 167 785 169 787
rect 103 767 105 772
rect 113 770 115 772
rect 148 775 150 777
rect 158 775 160 779
rect 167 776 169 782
rect 196 789 198 791
rect 201 789 204 791
rect 212 785 214 787
rect 148 767 150 772
rect 158 770 160 772
rect 193 775 195 777
rect 203 775 205 779
rect 212 776 214 782
rect 241 789 243 791
rect 246 789 249 791
rect 257 785 259 787
rect 193 767 195 772
rect 203 770 205 772
rect 238 775 240 777
rect 248 775 250 779
rect 257 776 259 782
rect 286 789 288 791
rect 291 789 294 791
rect 302 785 304 787
rect 238 767 240 772
rect 248 770 250 772
rect 283 775 285 777
rect 293 775 295 779
rect 302 776 304 782
rect 331 789 333 791
rect 336 789 339 791
rect 347 785 349 787
rect 283 767 285 772
rect 293 770 295 772
rect 328 775 330 777
rect 338 775 340 779
rect 347 776 349 782
rect 376 789 378 791
rect 381 789 384 791
rect 392 785 394 787
rect 328 767 330 772
rect 338 770 340 772
rect 373 775 375 777
rect 383 775 385 779
rect 392 776 394 782
rect 421 789 423 791
rect 426 789 429 791
rect 437 785 439 787
rect 373 767 375 772
rect 383 770 385 772
rect 418 775 420 777
rect 428 775 430 779
rect 437 776 439 782
rect 466 789 468 791
rect 471 789 474 791
rect 482 785 484 787
rect 418 767 420 772
rect 428 770 430 772
rect 463 775 465 777
rect 473 775 475 779
rect 482 776 484 782
rect 511 789 513 791
rect 516 789 519 791
rect 527 785 529 787
rect 463 767 465 772
rect 473 770 475 772
rect 508 775 510 777
rect 518 775 520 779
rect 527 776 529 782
rect 556 789 558 791
rect 561 789 564 791
rect 572 785 574 787
rect 508 767 510 772
rect 518 770 520 772
rect 553 775 555 777
rect 563 775 565 779
rect 572 776 574 782
rect 601 789 603 791
rect 606 789 609 791
rect 617 785 619 787
rect 553 767 555 772
rect 563 770 565 772
rect 598 775 600 777
rect 608 775 610 779
rect 617 776 619 782
rect 646 789 648 791
rect 651 789 654 791
rect 662 785 664 787
rect 598 767 600 772
rect 608 770 610 772
rect 643 775 645 777
rect 653 775 655 779
rect 662 776 664 782
rect 691 789 693 791
rect 696 789 699 791
rect 707 785 709 787
rect 643 767 645 772
rect 653 770 655 772
rect 688 775 690 777
rect 698 775 700 779
rect 707 776 709 782
rect 736 789 738 791
rect 741 789 744 791
rect 752 785 754 787
rect 688 767 690 772
rect 698 770 700 772
rect 733 775 735 777
rect 743 775 745 779
rect 752 776 754 782
rect 781 789 783 791
rect 786 789 789 791
rect 797 785 799 787
rect 733 767 735 772
rect 743 770 745 772
rect 778 775 780 777
rect 788 775 790 779
rect 797 776 799 782
rect 826 789 828 791
rect 831 789 834 791
rect 842 785 844 787
rect 778 767 780 772
rect 788 770 790 772
rect 823 775 825 777
rect 833 775 835 779
rect 842 776 844 782
rect 871 789 873 791
rect 876 789 879 791
rect 887 785 889 787
rect 823 767 825 772
rect 833 770 835 772
rect 868 775 870 777
rect 878 775 880 779
rect 887 776 889 782
rect 868 767 870 772
rect 878 770 880 772
rect 16 744 18 746
rect 21 744 24 746
rect 32 740 34 742
rect 13 730 15 732
rect 23 730 25 734
rect 32 731 34 737
rect 61 744 63 746
rect 66 744 69 746
rect 77 740 79 742
rect 13 722 15 727
rect 23 725 25 727
rect 58 730 60 732
rect 68 730 70 734
rect 77 731 79 737
rect 106 744 108 746
rect 111 744 114 746
rect 122 740 124 742
rect 58 722 60 727
rect 68 725 70 727
rect 103 730 105 732
rect 113 730 115 734
rect 122 731 124 737
rect 151 744 153 746
rect 156 744 159 746
rect 167 740 169 742
rect 103 722 105 727
rect 113 725 115 727
rect 148 730 150 732
rect 158 730 160 734
rect 167 731 169 737
rect 196 744 198 746
rect 201 744 204 746
rect 212 740 214 742
rect 148 722 150 727
rect 158 725 160 727
rect 193 730 195 732
rect 203 730 205 734
rect 212 731 214 737
rect 241 744 243 746
rect 246 744 249 746
rect 257 740 259 742
rect 193 722 195 727
rect 203 725 205 727
rect 238 730 240 732
rect 248 730 250 734
rect 257 731 259 737
rect 286 744 288 746
rect 291 744 294 746
rect 302 740 304 742
rect 238 722 240 727
rect 248 725 250 727
rect 283 730 285 732
rect 293 730 295 734
rect 302 731 304 737
rect 331 744 333 746
rect 336 744 339 746
rect 347 740 349 742
rect 283 722 285 727
rect 293 725 295 727
rect 328 730 330 732
rect 338 730 340 734
rect 347 731 349 737
rect 376 744 378 746
rect 381 744 384 746
rect 392 740 394 742
rect 328 722 330 727
rect 338 725 340 727
rect 373 730 375 732
rect 383 730 385 734
rect 392 731 394 737
rect 421 744 423 746
rect 426 744 429 746
rect 437 740 439 742
rect 373 722 375 727
rect 383 725 385 727
rect 418 730 420 732
rect 428 730 430 734
rect 437 731 439 737
rect 466 744 468 746
rect 471 744 474 746
rect 482 740 484 742
rect 418 722 420 727
rect 428 725 430 727
rect 463 730 465 732
rect 473 730 475 734
rect 482 731 484 737
rect 511 744 513 746
rect 516 744 519 746
rect 527 740 529 742
rect 463 722 465 727
rect 473 725 475 727
rect 508 730 510 732
rect 518 730 520 734
rect 527 731 529 737
rect 556 744 558 746
rect 561 744 564 746
rect 572 740 574 742
rect 508 722 510 727
rect 518 725 520 727
rect 553 730 555 732
rect 563 730 565 734
rect 572 731 574 737
rect 601 744 603 746
rect 606 744 609 746
rect 617 740 619 742
rect 553 722 555 727
rect 563 725 565 727
rect 598 730 600 732
rect 608 730 610 734
rect 617 731 619 737
rect 646 744 648 746
rect 651 744 654 746
rect 662 740 664 742
rect 598 722 600 727
rect 608 725 610 727
rect 643 730 645 732
rect 653 730 655 734
rect 662 731 664 737
rect 691 744 693 746
rect 696 744 699 746
rect 707 740 709 742
rect 643 722 645 727
rect 653 725 655 727
rect 688 730 690 732
rect 698 730 700 734
rect 707 731 709 737
rect 736 744 738 746
rect 741 744 744 746
rect 752 740 754 742
rect 688 722 690 727
rect 698 725 700 727
rect 733 730 735 732
rect 743 730 745 734
rect 752 731 754 737
rect 781 744 783 746
rect 786 744 789 746
rect 797 740 799 742
rect 733 722 735 727
rect 743 725 745 727
rect 778 730 780 732
rect 788 730 790 734
rect 797 731 799 737
rect 826 744 828 746
rect 831 744 834 746
rect 842 740 844 742
rect 778 722 780 727
rect 788 725 790 727
rect 823 730 825 732
rect 833 730 835 734
rect 842 731 844 737
rect 871 744 873 746
rect 876 744 879 746
rect 887 740 889 742
rect 823 722 825 727
rect 833 725 835 727
rect 868 730 870 732
rect 878 730 880 734
rect 887 731 889 737
rect 868 722 870 727
rect 878 725 880 727
rect 16 699 18 701
rect 21 699 24 701
rect 32 695 34 697
rect 13 685 15 687
rect 23 685 25 689
rect 32 686 34 692
rect 61 699 63 701
rect 66 699 69 701
rect 77 695 79 697
rect 13 677 15 682
rect 23 680 25 682
rect 58 685 60 687
rect 68 685 70 689
rect 77 686 79 692
rect 106 699 108 701
rect 111 699 114 701
rect 122 695 124 697
rect 58 677 60 682
rect 68 680 70 682
rect 103 685 105 687
rect 113 685 115 689
rect 122 686 124 692
rect 151 699 153 701
rect 156 699 159 701
rect 167 695 169 697
rect 103 677 105 682
rect 113 680 115 682
rect 148 685 150 687
rect 158 685 160 689
rect 167 686 169 692
rect 196 699 198 701
rect 201 699 204 701
rect 212 695 214 697
rect 148 677 150 682
rect 158 680 160 682
rect 193 685 195 687
rect 203 685 205 689
rect 212 686 214 692
rect 241 699 243 701
rect 246 699 249 701
rect 257 695 259 697
rect 193 677 195 682
rect 203 680 205 682
rect 238 685 240 687
rect 248 685 250 689
rect 257 686 259 692
rect 286 699 288 701
rect 291 699 294 701
rect 302 695 304 697
rect 238 677 240 682
rect 248 680 250 682
rect 283 685 285 687
rect 293 685 295 689
rect 302 686 304 692
rect 331 699 333 701
rect 336 699 339 701
rect 347 695 349 697
rect 283 677 285 682
rect 293 680 295 682
rect 328 685 330 687
rect 338 685 340 689
rect 347 686 349 692
rect 376 699 378 701
rect 381 699 384 701
rect 392 695 394 697
rect 328 677 330 682
rect 338 680 340 682
rect 373 685 375 687
rect 383 685 385 689
rect 392 686 394 692
rect 421 699 423 701
rect 426 699 429 701
rect 437 695 439 697
rect 373 677 375 682
rect 383 680 385 682
rect 418 685 420 687
rect 428 685 430 689
rect 437 686 439 692
rect 466 699 468 701
rect 471 699 474 701
rect 482 695 484 697
rect 418 677 420 682
rect 428 680 430 682
rect 463 685 465 687
rect 473 685 475 689
rect 482 686 484 692
rect 511 699 513 701
rect 516 699 519 701
rect 527 695 529 697
rect 463 677 465 682
rect 473 680 475 682
rect 508 685 510 687
rect 518 685 520 689
rect 527 686 529 692
rect 556 699 558 701
rect 561 699 564 701
rect 572 695 574 697
rect 508 677 510 682
rect 518 680 520 682
rect 553 685 555 687
rect 563 685 565 689
rect 572 686 574 692
rect 601 699 603 701
rect 606 699 609 701
rect 617 695 619 697
rect 553 677 555 682
rect 563 680 565 682
rect 598 685 600 687
rect 608 685 610 689
rect 617 686 619 692
rect 646 699 648 701
rect 651 699 654 701
rect 662 695 664 697
rect 598 677 600 682
rect 608 680 610 682
rect 643 685 645 687
rect 653 685 655 689
rect 662 686 664 692
rect 691 699 693 701
rect 696 699 699 701
rect 707 695 709 697
rect 643 677 645 682
rect 653 680 655 682
rect 688 685 690 687
rect 698 685 700 689
rect 707 686 709 692
rect 736 699 738 701
rect 741 699 744 701
rect 752 695 754 697
rect 688 677 690 682
rect 698 680 700 682
rect 733 685 735 687
rect 743 685 745 689
rect 752 686 754 692
rect 781 699 783 701
rect 786 699 789 701
rect 797 695 799 697
rect 733 677 735 682
rect 743 680 745 682
rect 778 685 780 687
rect 788 685 790 689
rect 797 686 799 692
rect 826 699 828 701
rect 831 699 834 701
rect 842 695 844 697
rect 778 677 780 682
rect 788 680 790 682
rect 823 685 825 687
rect 833 685 835 689
rect 842 686 844 692
rect 871 699 873 701
rect 876 699 879 701
rect 887 695 889 697
rect 823 677 825 682
rect 833 680 835 682
rect 868 685 870 687
rect 878 685 880 689
rect 887 686 889 692
rect 868 677 870 682
rect 878 680 880 682
rect 16 654 18 656
rect 21 654 24 656
rect 32 650 34 652
rect 13 640 15 642
rect 23 640 25 644
rect 32 641 34 647
rect 61 654 63 656
rect 66 654 69 656
rect 77 650 79 652
rect 13 632 15 637
rect 23 635 25 637
rect 58 640 60 642
rect 68 640 70 644
rect 77 641 79 647
rect 106 654 108 656
rect 111 654 114 656
rect 122 650 124 652
rect 58 632 60 637
rect 68 635 70 637
rect 103 640 105 642
rect 113 640 115 644
rect 122 641 124 647
rect 151 654 153 656
rect 156 654 159 656
rect 167 650 169 652
rect 103 632 105 637
rect 113 635 115 637
rect 148 640 150 642
rect 158 640 160 644
rect 167 641 169 647
rect 196 654 198 656
rect 201 654 204 656
rect 212 650 214 652
rect 148 632 150 637
rect 158 635 160 637
rect 193 640 195 642
rect 203 640 205 644
rect 212 641 214 647
rect 241 654 243 656
rect 246 654 249 656
rect 257 650 259 652
rect 193 632 195 637
rect 203 635 205 637
rect 238 640 240 642
rect 248 640 250 644
rect 257 641 259 647
rect 286 654 288 656
rect 291 654 294 656
rect 302 650 304 652
rect 238 632 240 637
rect 248 635 250 637
rect 283 640 285 642
rect 293 640 295 644
rect 302 641 304 647
rect 331 654 333 656
rect 336 654 339 656
rect 347 650 349 652
rect 283 632 285 637
rect 293 635 295 637
rect 328 640 330 642
rect 338 640 340 644
rect 347 641 349 647
rect 376 654 378 656
rect 381 654 384 656
rect 392 650 394 652
rect 328 632 330 637
rect 338 635 340 637
rect 373 640 375 642
rect 383 640 385 644
rect 392 641 394 647
rect 421 654 423 656
rect 426 654 429 656
rect 437 650 439 652
rect 373 632 375 637
rect 383 635 385 637
rect 418 640 420 642
rect 428 640 430 644
rect 437 641 439 647
rect 466 654 468 656
rect 471 654 474 656
rect 482 650 484 652
rect 418 632 420 637
rect 428 635 430 637
rect 463 640 465 642
rect 473 640 475 644
rect 482 641 484 647
rect 511 654 513 656
rect 516 654 519 656
rect 527 650 529 652
rect 463 632 465 637
rect 473 635 475 637
rect 508 640 510 642
rect 518 640 520 644
rect 527 641 529 647
rect 556 654 558 656
rect 561 654 564 656
rect 572 650 574 652
rect 508 632 510 637
rect 518 635 520 637
rect 553 640 555 642
rect 563 640 565 644
rect 572 641 574 647
rect 601 654 603 656
rect 606 654 609 656
rect 617 650 619 652
rect 553 632 555 637
rect 563 635 565 637
rect 598 640 600 642
rect 608 640 610 644
rect 617 641 619 647
rect 646 654 648 656
rect 651 654 654 656
rect 662 650 664 652
rect 598 632 600 637
rect 608 635 610 637
rect 643 640 645 642
rect 653 640 655 644
rect 662 641 664 647
rect 691 654 693 656
rect 696 654 699 656
rect 707 650 709 652
rect 643 632 645 637
rect 653 635 655 637
rect 688 640 690 642
rect 698 640 700 644
rect 707 641 709 647
rect 736 654 738 656
rect 741 654 744 656
rect 752 650 754 652
rect 688 632 690 637
rect 698 635 700 637
rect 733 640 735 642
rect 743 640 745 644
rect 752 641 754 647
rect 781 654 783 656
rect 786 654 789 656
rect 797 650 799 652
rect 733 632 735 637
rect 743 635 745 637
rect 778 640 780 642
rect 788 640 790 644
rect 797 641 799 647
rect 826 654 828 656
rect 831 654 834 656
rect 842 650 844 652
rect 778 632 780 637
rect 788 635 790 637
rect 823 640 825 642
rect 833 640 835 644
rect 842 641 844 647
rect 871 654 873 656
rect 876 654 879 656
rect 887 650 889 652
rect 823 632 825 637
rect 833 635 835 637
rect 868 640 870 642
rect 878 640 880 644
rect 887 641 889 647
rect 868 632 870 637
rect 878 635 880 637
rect 16 609 18 611
rect 21 609 24 611
rect 32 605 34 607
rect 13 595 15 597
rect 23 595 25 599
rect 32 596 34 602
rect 61 609 63 611
rect 66 609 69 611
rect 77 605 79 607
rect 13 587 15 592
rect 23 590 25 592
rect 58 595 60 597
rect 68 595 70 599
rect 77 596 79 602
rect 106 609 108 611
rect 111 609 114 611
rect 122 605 124 607
rect 58 587 60 592
rect 68 590 70 592
rect 103 595 105 597
rect 113 595 115 599
rect 122 596 124 602
rect 151 609 153 611
rect 156 609 159 611
rect 167 605 169 607
rect 103 587 105 592
rect 113 590 115 592
rect 148 595 150 597
rect 158 595 160 599
rect 167 596 169 602
rect 196 609 198 611
rect 201 609 204 611
rect 212 605 214 607
rect 148 587 150 592
rect 158 590 160 592
rect 193 595 195 597
rect 203 595 205 599
rect 212 596 214 602
rect 241 609 243 611
rect 246 609 249 611
rect 257 605 259 607
rect 193 587 195 592
rect 203 590 205 592
rect 238 595 240 597
rect 248 595 250 599
rect 257 596 259 602
rect 286 609 288 611
rect 291 609 294 611
rect 302 605 304 607
rect 238 587 240 592
rect 248 590 250 592
rect 283 595 285 597
rect 293 595 295 599
rect 302 596 304 602
rect 331 609 333 611
rect 336 609 339 611
rect 347 605 349 607
rect 283 587 285 592
rect 293 590 295 592
rect 328 595 330 597
rect 338 595 340 599
rect 347 596 349 602
rect 376 609 378 611
rect 381 609 384 611
rect 392 605 394 607
rect 328 587 330 592
rect 338 590 340 592
rect 373 595 375 597
rect 383 595 385 599
rect 392 596 394 602
rect 421 609 423 611
rect 426 609 429 611
rect 437 605 439 607
rect 373 587 375 592
rect 383 590 385 592
rect 418 595 420 597
rect 428 595 430 599
rect 437 596 439 602
rect 466 609 468 611
rect 471 609 474 611
rect 482 605 484 607
rect 418 587 420 592
rect 428 590 430 592
rect 463 595 465 597
rect 473 595 475 599
rect 482 596 484 602
rect 511 609 513 611
rect 516 609 519 611
rect 527 605 529 607
rect 463 587 465 592
rect 473 590 475 592
rect 508 595 510 597
rect 518 595 520 599
rect 527 596 529 602
rect 556 609 558 611
rect 561 609 564 611
rect 572 605 574 607
rect 508 587 510 592
rect 518 590 520 592
rect 553 595 555 597
rect 563 595 565 599
rect 572 596 574 602
rect 601 609 603 611
rect 606 609 609 611
rect 617 605 619 607
rect 553 587 555 592
rect 563 590 565 592
rect 598 595 600 597
rect 608 595 610 599
rect 617 596 619 602
rect 646 609 648 611
rect 651 609 654 611
rect 662 605 664 607
rect 598 587 600 592
rect 608 590 610 592
rect 643 595 645 597
rect 653 595 655 599
rect 662 596 664 602
rect 691 609 693 611
rect 696 609 699 611
rect 707 605 709 607
rect 643 587 645 592
rect 653 590 655 592
rect 688 595 690 597
rect 698 595 700 599
rect 707 596 709 602
rect 736 609 738 611
rect 741 609 744 611
rect 752 605 754 607
rect 688 587 690 592
rect 698 590 700 592
rect 733 595 735 597
rect 743 595 745 599
rect 752 596 754 602
rect 781 609 783 611
rect 786 609 789 611
rect 797 605 799 607
rect 733 587 735 592
rect 743 590 745 592
rect 778 595 780 597
rect 788 595 790 599
rect 797 596 799 602
rect 826 609 828 611
rect 831 609 834 611
rect 842 605 844 607
rect 778 587 780 592
rect 788 590 790 592
rect 823 595 825 597
rect 833 595 835 599
rect 842 596 844 602
rect 871 609 873 611
rect 876 609 879 611
rect 887 605 889 607
rect 823 587 825 592
rect 833 590 835 592
rect 868 595 870 597
rect 878 595 880 599
rect 887 596 889 602
rect 868 587 870 592
rect 878 590 880 592
rect 16 564 18 566
rect 21 564 24 566
rect 32 560 34 562
rect 13 550 15 552
rect 23 550 25 554
rect 32 551 34 557
rect 61 564 63 566
rect 66 564 69 566
rect 77 560 79 562
rect 13 542 15 547
rect 23 545 25 547
rect 58 550 60 552
rect 68 550 70 554
rect 77 551 79 557
rect 106 564 108 566
rect 111 564 114 566
rect 122 560 124 562
rect 58 542 60 547
rect 68 545 70 547
rect 103 550 105 552
rect 113 550 115 554
rect 122 551 124 557
rect 151 564 153 566
rect 156 564 159 566
rect 167 560 169 562
rect 103 542 105 547
rect 113 545 115 547
rect 148 550 150 552
rect 158 550 160 554
rect 167 551 169 557
rect 196 564 198 566
rect 201 564 204 566
rect 212 560 214 562
rect 148 542 150 547
rect 158 545 160 547
rect 193 550 195 552
rect 203 550 205 554
rect 212 551 214 557
rect 241 564 243 566
rect 246 564 249 566
rect 257 560 259 562
rect 193 542 195 547
rect 203 545 205 547
rect 238 550 240 552
rect 248 550 250 554
rect 257 551 259 557
rect 286 564 288 566
rect 291 564 294 566
rect 302 560 304 562
rect 238 542 240 547
rect 248 545 250 547
rect 283 550 285 552
rect 293 550 295 554
rect 302 551 304 557
rect 331 564 333 566
rect 336 564 339 566
rect 347 560 349 562
rect 283 542 285 547
rect 293 545 295 547
rect 328 550 330 552
rect 338 550 340 554
rect 347 551 349 557
rect 376 564 378 566
rect 381 564 384 566
rect 392 560 394 562
rect 328 542 330 547
rect 338 545 340 547
rect 373 550 375 552
rect 383 550 385 554
rect 392 551 394 557
rect 421 564 423 566
rect 426 564 429 566
rect 437 560 439 562
rect 373 542 375 547
rect 383 545 385 547
rect 418 550 420 552
rect 428 550 430 554
rect 437 551 439 557
rect 466 564 468 566
rect 471 564 474 566
rect 482 560 484 562
rect 418 542 420 547
rect 428 545 430 547
rect 463 550 465 552
rect 473 550 475 554
rect 482 551 484 557
rect 511 564 513 566
rect 516 564 519 566
rect 527 560 529 562
rect 463 542 465 547
rect 473 545 475 547
rect 508 550 510 552
rect 518 550 520 554
rect 527 551 529 557
rect 556 564 558 566
rect 561 564 564 566
rect 572 560 574 562
rect 508 542 510 547
rect 518 545 520 547
rect 553 550 555 552
rect 563 550 565 554
rect 572 551 574 557
rect 601 564 603 566
rect 606 564 609 566
rect 617 560 619 562
rect 553 542 555 547
rect 563 545 565 547
rect 598 550 600 552
rect 608 550 610 554
rect 617 551 619 557
rect 646 564 648 566
rect 651 564 654 566
rect 662 560 664 562
rect 598 542 600 547
rect 608 545 610 547
rect 643 550 645 552
rect 653 550 655 554
rect 662 551 664 557
rect 691 564 693 566
rect 696 564 699 566
rect 707 560 709 562
rect 643 542 645 547
rect 653 545 655 547
rect 688 550 690 552
rect 698 550 700 554
rect 707 551 709 557
rect 736 564 738 566
rect 741 564 744 566
rect 752 560 754 562
rect 688 542 690 547
rect 698 545 700 547
rect 733 550 735 552
rect 743 550 745 554
rect 752 551 754 557
rect 781 564 783 566
rect 786 564 789 566
rect 797 560 799 562
rect 733 542 735 547
rect 743 545 745 547
rect 778 550 780 552
rect 788 550 790 554
rect 797 551 799 557
rect 826 564 828 566
rect 831 564 834 566
rect 842 560 844 562
rect 778 542 780 547
rect 788 545 790 547
rect 823 550 825 552
rect 833 550 835 554
rect 842 551 844 557
rect 871 564 873 566
rect 876 564 879 566
rect 887 560 889 562
rect 823 542 825 547
rect 833 545 835 547
rect 868 550 870 552
rect 878 550 880 554
rect 887 551 889 557
rect 868 542 870 547
rect 878 545 880 547
rect 16 519 18 521
rect 21 519 24 521
rect 32 515 34 517
rect 13 505 15 507
rect 23 505 25 509
rect 32 506 34 512
rect 61 519 63 521
rect 66 519 69 521
rect 77 515 79 517
rect 13 497 15 502
rect 23 500 25 502
rect 58 505 60 507
rect 68 505 70 509
rect 77 506 79 512
rect 106 519 108 521
rect 111 519 114 521
rect 122 515 124 517
rect 58 497 60 502
rect 68 500 70 502
rect 103 505 105 507
rect 113 505 115 509
rect 122 506 124 512
rect 151 519 153 521
rect 156 519 159 521
rect 167 515 169 517
rect 103 497 105 502
rect 113 500 115 502
rect 148 505 150 507
rect 158 505 160 509
rect 167 506 169 512
rect 196 519 198 521
rect 201 519 204 521
rect 212 515 214 517
rect 148 497 150 502
rect 158 500 160 502
rect 193 505 195 507
rect 203 505 205 509
rect 212 506 214 512
rect 241 519 243 521
rect 246 519 249 521
rect 257 515 259 517
rect 193 497 195 502
rect 203 500 205 502
rect 238 505 240 507
rect 248 505 250 509
rect 257 506 259 512
rect 286 519 288 521
rect 291 519 294 521
rect 302 515 304 517
rect 238 497 240 502
rect 248 500 250 502
rect 283 505 285 507
rect 293 505 295 509
rect 302 506 304 512
rect 331 519 333 521
rect 336 519 339 521
rect 347 515 349 517
rect 283 497 285 502
rect 293 500 295 502
rect 328 505 330 507
rect 338 505 340 509
rect 347 506 349 512
rect 376 519 378 521
rect 381 519 384 521
rect 392 515 394 517
rect 328 497 330 502
rect 338 500 340 502
rect 373 505 375 507
rect 383 505 385 509
rect 392 506 394 512
rect 421 519 423 521
rect 426 519 429 521
rect 437 515 439 517
rect 373 497 375 502
rect 383 500 385 502
rect 418 505 420 507
rect 428 505 430 509
rect 437 506 439 512
rect 466 519 468 521
rect 471 519 474 521
rect 482 515 484 517
rect 418 497 420 502
rect 428 500 430 502
rect 463 505 465 507
rect 473 505 475 509
rect 482 506 484 512
rect 511 519 513 521
rect 516 519 519 521
rect 527 515 529 517
rect 463 497 465 502
rect 473 500 475 502
rect 508 505 510 507
rect 518 505 520 509
rect 527 506 529 512
rect 556 519 558 521
rect 561 519 564 521
rect 572 515 574 517
rect 508 497 510 502
rect 518 500 520 502
rect 553 505 555 507
rect 563 505 565 509
rect 572 506 574 512
rect 601 519 603 521
rect 606 519 609 521
rect 617 515 619 517
rect 553 497 555 502
rect 563 500 565 502
rect 598 505 600 507
rect 608 505 610 509
rect 617 506 619 512
rect 646 519 648 521
rect 651 519 654 521
rect 662 515 664 517
rect 598 497 600 502
rect 608 500 610 502
rect 643 505 645 507
rect 653 505 655 509
rect 662 506 664 512
rect 691 519 693 521
rect 696 519 699 521
rect 707 515 709 517
rect 643 497 645 502
rect 653 500 655 502
rect 688 505 690 507
rect 698 505 700 509
rect 707 506 709 512
rect 736 519 738 521
rect 741 519 744 521
rect 752 515 754 517
rect 688 497 690 502
rect 698 500 700 502
rect 733 505 735 507
rect 743 505 745 509
rect 752 506 754 512
rect 781 519 783 521
rect 786 519 789 521
rect 797 515 799 517
rect 733 497 735 502
rect 743 500 745 502
rect 778 505 780 507
rect 788 505 790 509
rect 797 506 799 512
rect 826 519 828 521
rect 831 519 834 521
rect 842 515 844 517
rect 778 497 780 502
rect 788 500 790 502
rect 823 505 825 507
rect 833 505 835 509
rect 842 506 844 512
rect 871 519 873 521
rect 876 519 879 521
rect 887 515 889 517
rect 823 497 825 502
rect 833 500 835 502
rect 868 505 870 507
rect 878 505 880 509
rect 887 506 889 512
rect 868 497 870 502
rect 878 500 880 502
rect 16 474 18 476
rect 21 474 24 476
rect 32 470 34 472
rect 13 460 15 462
rect 23 460 25 464
rect 32 461 34 467
rect 61 474 63 476
rect 66 474 69 476
rect 77 470 79 472
rect 13 452 15 457
rect 23 455 25 457
rect 58 460 60 462
rect 68 460 70 464
rect 77 461 79 467
rect 106 474 108 476
rect 111 474 114 476
rect 122 470 124 472
rect 58 452 60 457
rect 68 455 70 457
rect 103 460 105 462
rect 113 460 115 464
rect 122 461 124 467
rect 151 474 153 476
rect 156 474 159 476
rect 167 470 169 472
rect 103 452 105 457
rect 113 455 115 457
rect 148 460 150 462
rect 158 460 160 464
rect 167 461 169 467
rect 196 474 198 476
rect 201 474 204 476
rect 212 470 214 472
rect 148 452 150 457
rect 158 455 160 457
rect 193 460 195 462
rect 203 460 205 464
rect 212 461 214 467
rect 241 474 243 476
rect 246 474 249 476
rect 257 470 259 472
rect 193 452 195 457
rect 203 455 205 457
rect 238 460 240 462
rect 248 460 250 464
rect 257 461 259 467
rect 286 474 288 476
rect 291 474 294 476
rect 302 470 304 472
rect 238 452 240 457
rect 248 455 250 457
rect 283 460 285 462
rect 293 460 295 464
rect 302 461 304 467
rect 331 474 333 476
rect 336 474 339 476
rect 347 470 349 472
rect 283 452 285 457
rect 293 455 295 457
rect 328 460 330 462
rect 338 460 340 464
rect 347 461 349 467
rect 376 474 378 476
rect 381 474 384 476
rect 392 470 394 472
rect 328 452 330 457
rect 338 455 340 457
rect 373 460 375 462
rect 383 460 385 464
rect 392 461 394 467
rect 421 474 423 476
rect 426 474 429 476
rect 437 470 439 472
rect 373 452 375 457
rect 383 455 385 457
rect 418 460 420 462
rect 428 460 430 464
rect 437 461 439 467
rect 466 474 468 476
rect 471 474 474 476
rect 482 470 484 472
rect 418 452 420 457
rect 428 455 430 457
rect 463 460 465 462
rect 473 460 475 464
rect 482 461 484 467
rect 511 474 513 476
rect 516 474 519 476
rect 527 470 529 472
rect 463 452 465 457
rect 473 455 475 457
rect 508 460 510 462
rect 518 460 520 464
rect 527 461 529 467
rect 556 474 558 476
rect 561 474 564 476
rect 572 470 574 472
rect 508 452 510 457
rect 518 455 520 457
rect 553 460 555 462
rect 563 460 565 464
rect 572 461 574 467
rect 601 474 603 476
rect 606 474 609 476
rect 617 470 619 472
rect 553 452 555 457
rect 563 455 565 457
rect 598 460 600 462
rect 608 460 610 464
rect 617 461 619 467
rect 646 474 648 476
rect 651 474 654 476
rect 662 470 664 472
rect 598 452 600 457
rect 608 455 610 457
rect 643 460 645 462
rect 653 460 655 464
rect 662 461 664 467
rect 691 474 693 476
rect 696 474 699 476
rect 707 470 709 472
rect 643 452 645 457
rect 653 455 655 457
rect 688 460 690 462
rect 698 460 700 464
rect 707 461 709 467
rect 736 474 738 476
rect 741 474 744 476
rect 752 470 754 472
rect 688 452 690 457
rect 698 455 700 457
rect 733 460 735 462
rect 743 460 745 464
rect 752 461 754 467
rect 781 474 783 476
rect 786 474 789 476
rect 797 470 799 472
rect 733 452 735 457
rect 743 455 745 457
rect 778 460 780 462
rect 788 460 790 464
rect 797 461 799 467
rect 826 474 828 476
rect 831 474 834 476
rect 842 470 844 472
rect 778 452 780 457
rect 788 455 790 457
rect 823 460 825 462
rect 833 460 835 464
rect 842 461 844 467
rect 871 474 873 476
rect 876 474 879 476
rect 887 470 889 472
rect 823 452 825 457
rect 833 455 835 457
rect 868 460 870 462
rect 878 460 880 464
rect 887 461 889 467
rect 868 452 870 457
rect 878 455 880 457
rect 16 429 18 431
rect 21 429 24 431
rect 32 425 34 427
rect 13 415 15 417
rect 23 415 25 419
rect 32 416 34 422
rect 61 429 63 431
rect 66 429 69 431
rect 77 425 79 427
rect 13 407 15 412
rect 23 410 25 412
rect 58 415 60 417
rect 68 415 70 419
rect 77 416 79 422
rect 106 429 108 431
rect 111 429 114 431
rect 122 425 124 427
rect 58 407 60 412
rect 68 410 70 412
rect 103 415 105 417
rect 113 415 115 419
rect 122 416 124 422
rect 151 429 153 431
rect 156 429 159 431
rect 167 425 169 427
rect 103 407 105 412
rect 113 410 115 412
rect 148 415 150 417
rect 158 415 160 419
rect 167 416 169 422
rect 196 429 198 431
rect 201 429 204 431
rect 212 425 214 427
rect 148 407 150 412
rect 158 410 160 412
rect 193 415 195 417
rect 203 415 205 419
rect 212 416 214 422
rect 241 429 243 431
rect 246 429 249 431
rect 257 425 259 427
rect 193 407 195 412
rect 203 410 205 412
rect 238 415 240 417
rect 248 415 250 419
rect 257 416 259 422
rect 286 429 288 431
rect 291 429 294 431
rect 302 425 304 427
rect 238 407 240 412
rect 248 410 250 412
rect 283 415 285 417
rect 293 415 295 419
rect 302 416 304 422
rect 331 429 333 431
rect 336 429 339 431
rect 347 425 349 427
rect 283 407 285 412
rect 293 410 295 412
rect 328 415 330 417
rect 338 415 340 419
rect 347 416 349 422
rect 376 429 378 431
rect 381 429 384 431
rect 392 425 394 427
rect 328 407 330 412
rect 338 410 340 412
rect 373 415 375 417
rect 383 415 385 419
rect 392 416 394 422
rect 421 429 423 431
rect 426 429 429 431
rect 437 425 439 427
rect 373 407 375 412
rect 383 410 385 412
rect 418 415 420 417
rect 428 415 430 419
rect 437 416 439 422
rect 466 429 468 431
rect 471 429 474 431
rect 482 425 484 427
rect 418 407 420 412
rect 428 410 430 412
rect 463 415 465 417
rect 473 415 475 419
rect 482 416 484 422
rect 511 429 513 431
rect 516 429 519 431
rect 527 425 529 427
rect 463 407 465 412
rect 473 410 475 412
rect 508 415 510 417
rect 518 415 520 419
rect 527 416 529 422
rect 556 429 558 431
rect 561 429 564 431
rect 572 425 574 427
rect 508 407 510 412
rect 518 410 520 412
rect 553 415 555 417
rect 563 415 565 419
rect 572 416 574 422
rect 601 429 603 431
rect 606 429 609 431
rect 617 425 619 427
rect 553 407 555 412
rect 563 410 565 412
rect 598 415 600 417
rect 608 415 610 419
rect 617 416 619 422
rect 646 429 648 431
rect 651 429 654 431
rect 662 425 664 427
rect 598 407 600 412
rect 608 410 610 412
rect 643 415 645 417
rect 653 415 655 419
rect 662 416 664 422
rect 691 429 693 431
rect 696 429 699 431
rect 707 425 709 427
rect 643 407 645 412
rect 653 410 655 412
rect 688 415 690 417
rect 698 415 700 419
rect 707 416 709 422
rect 736 429 738 431
rect 741 429 744 431
rect 752 425 754 427
rect 688 407 690 412
rect 698 410 700 412
rect 733 415 735 417
rect 743 415 745 419
rect 752 416 754 422
rect 781 429 783 431
rect 786 429 789 431
rect 797 425 799 427
rect 733 407 735 412
rect 743 410 745 412
rect 778 415 780 417
rect 788 415 790 419
rect 797 416 799 422
rect 826 429 828 431
rect 831 429 834 431
rect 842 425 844 427
rect 778 407 780 412
rect 788 410 790 412
rect 823 415 825 417
rect 833 415 835 419
rect 842 416 844 422
rect 871 429 873 431
rect 876 429 879 431
rect 887 425 889 427
rect 823 407 825 412
rect 833 410 835 412
rect 868 415 870 417
rect 878 415 880 419
rect 887 416 889 422
rect 868 407 870 412
rect 878 410 880 412
rect 16 384 18 386
rect 21 384 24 386
rect 32 380 34 382
rect 13 370 15 372
rect 23 370 25 374
rect 32 371 34 377
rect 61 384 63 386
rect 66 384 69 386
rect 77 380 79 382
rect 13 362 15 367
rect 23 365 25 367
rect 58 370 60 372
rect 68 370 70 374
rect 77 371 79 377
rect 106 384 108 386
rect 111 384 114 386
rect 122 380 124 382
rect 58 362 60 367
rect 68 365 70 367
rect 103 370 105 372
rect 113 370 115 374
rect 122 371 124 377
rect 151 384 153 386
rect 156 384 159 386
rect 167 380 169 382
rect 103 362 105 367
rect 113 365 115 367
rect 148 370 150 372
rect 158 370 160 374
rect 167 371 169 377
rect 196 384 198 386
rect 201 384 204 386
rect 212 380 214 382
rect 148 362 150 367
rect 158 365 160 367
rect 193 370 195 372
rect 203 370 205 374
rect 212 371 214 377
rect 241 384 243 386
rect 246 384 249 386
rect 257 380 259 382
rect 193 362 195 367
rect 203 365 205 367
rect 238 370 240 372
rect 248 370 250 374
rect 257 371 259 377
rect 286 384 288 386
rect 291 384 294 386
rect 302 380 304 382
rect 238 362 240 367
rect 248 365 250 367
rect 283 370 285 372
rect 293 370 295 374
rect 302 371 304 377
rect 331 384 333 386
rect 336 384 339 386
rect 347 380 349 382
rect 283 362 285 367
rect 293 365 295 367
rect 328 370 330 372
rect 338 370 340 374
rect 347 371 349 377
rect 376 384 378 386
rect 381 384 384 386
rect 392 380 394 382
rect 328 362 330 367
rect 338 365 340 367
rect 373 370 375 372
rect 383 370 385 374
rect 392 371 394 377
rect 421 384 423 386
rect 426 384 429 386
rect 437 380 439 382
rect 373 362 375 367
rect 383 365 385 367
rect 418 370 420 372
rect 428 370 430 374
rect 437 371 439 377
rect 466 384 468 386
rect 471 384 474 386
rect 482 380 484 382
rect 418 362 420 367
rect 428 365 430 367
rect 463 370 465 372
rect 473 370 475 374
rect 482 371 484 377
rect 511 384 513 386
rect 516 384 519 386
rect 527 380 529 382
rect 463 362 465 367
rect 473 365 475 367
rect 508 370 510 372
rect 518 370 520 374
rect 527 371 529 377
rect 556 384 558 386
rect 561 384 564 386
rect 572 380 574 382
rect 508 362 510 367
rect 518 365 520 367
rect 553 370 555 372
rect 563 370 565 374
rect 572 371 574 377
rect 601 384 603 386
rect 606 384 609 386
rect 617 380 619 382
rect 553 362 555 367
rect 563 365 565 367
rect 598 370 600 372
rect 608 370 610 374
rect 617 371 619 377
rect 646 384 648 386
rect 651 384 654 386
rect 662 380 664 382
rect 598 362 600 367
rect 608 365 610 367
rect 643 370 645 372
rect 653 370 655 374
rect 662 371 664 377
rect 691 384 693 386
rect 696 384 699 386
rect 707 380 709 382
rect 643 362 645 367
rect 653 365 655 367
rect 688 370 690 372
rect 698 370 700 374
rect 707 371 709 377
rect 736 384 738 386
rect 741 384 744 386
rect 752 380 754 382
rect 688 362 690 367
rect 698 365 700 367
rect 733 370 735 372
rect 743 370 745 374
rect 752 371 754 377
rect 781 384 783 386
rect 786 384 789 386
rect 797 380 799 382
rect 733 362 735 367
rect 743 365 745 367
rect 778 370 780 372
rect 788 370 790 374
rect 797 371 799 377
rect 826 384 828 386
rect 831 384 834 386
rect 842 380 844 382
rect 778 362 780 367
rect 788 365 790 367
rect 823 370 825 372
rect 833 370 835 374
rect 842 371 844 377
rect 871 384 873 386
rect 876 384 879 386
rect 887 380 889 382
rect 823 362 825 367
rect 833 365 835 367
rect 868 370 870 372
rect 878 370 880 374
rect 887 371 889 377
rect 868 362 870 367
rect 878 365 880 367
rect 16 339 18 341
rect 21 339 24 341
rect 32 335 34 337
rect 13 325 15 327
rect 23 325 25 329
rect 32 326 34 332
rect 61 339 63 341
rect 66 339 69 341
rect 77 335 79 337
rect 13 317 15 322
rect 23 320 25 322
rect 58 325 60 327
rect 68 325 70 329
rect 77 326 79 332
rect 106 339 108 341
rect 111 339 114 341
rect 122 335 124 337
rect 58 317 60 322
rect 68 320 70 322
rect 103 325 105 327
rect 113 325 115 329
rect 122 326 124 332
rect 151 339 153 341
rect 156 339 159 341
rect 167 335 169 337
rect 103 317 105 322
rect 113 320 115 322
rect 148 325 150 327
rect 158 325 160 329
rect 167 326 169 332
rect 196 339 198 341
rect 201 339 204 341
rect 212 335 214 337
rect 148 317 150 322
rect 158 320 160 322
rect 193 325 195 327
rect 203 325 205 329
rect 212 326 214 332
rect 241 339 243 341
rect 246 339 249 341
rect 257 335 259 337
rect 193 317 195 322
rect 203 320 205 322
rect 238 325 240 327
rect 248 325 250 329
rect 257 326 259 332
rect 286 339 288 341
rect 291 339 294 341
rect 302 335 304 337
rect 238 317 240 322
rect 248 320 250 322
rect 283 325 285 327
rect 293 325 295 329
rect 302 326 304 332
rect 331 339 333 341
rect 336 339 339 341
rect 347 335 349 337
rect 283 317 285 322
rect 293 320 295 322
rect 328 325 330 327
rect 338 325 340 329
rect 347 326 349 332
rect 376 339 378 341
rect 381 339 384 341
rect 392 335 394 337
rect 328 317 330 322
rect 338 320 340 322
rect 373 325 375 327
rect 383 325 385 329
rect 392 326 394 332
rect 421 339 423 341
rect 426 339 429 341
rect 437 335 439 337
rect 373 317 375 322
rect 383 320 385 322
rect 418 325 420 327
rect 428 325 430 329
rect 437 326 439 332
rect 466 339 468 341
rect 471 339 474 341
rect 482 335 484 337
rect 418 317 420 322
rect 428 320 430 322
rect 463 325 465 327
rect 473 325 475 329
rect 482 326 484 332
rect 511 339 513 341
rect 516 339 519 341
rect 527 335 529 337
rect 463 317 465 322
rect 473 320 475 322
rect 508 325 510 327
rect 518 325 520 329
rect 527 326 529 332
rect 556 339 558 341
rect 561 339 564 341
rect 572 335 574 337
rect 508 317 510 322
rect 518 320 520 322
rect 553 325 555 327
rect 563 325 565 329
rect 572 326 574 332
rect 601 339 603 341
rect 606 339 609 341
rect 617 335 619 337
rect 553 317 555 322
rect 563 320 565 322
rect 598 325 600 327
rect 608 325 610 329
rect 617 326 619 332
rect 646 339 648 341
rect 651 339 654 341
rect 662 335 664 337
rect 598 317 600 322
rect 608 320 610 322
rect 643 325 645 327
rect 653 325 655 329
rect 662 326 664 332
rect 691 339 693 341
rect 696 339 699 341
rect 707 335 709 337
rect 643 317 645 322
rect 653 320 655 322
rect 688 325 690 327
rect 698 325 700 329
rect 707 326 709 332
rect 736 339 738 341
rect 741 339 744 341
rect 752 335 754 337
rect 688 317 690 322
rect 698 320 700 322
rect 733 325 735 327
rect 743 325 745 329
rect 752 326 754 332
rect 781 339 783 341
rect 786 339 789 341
rect 797 335 799 337
rect 733 317 735 322
rect 743 320 745 322
rect 778 325 780 327
rect 788 325 790 329
rect 797 326 799 332
rect 826 339 828 341
rect 831 339 834 341
rect 842 335 844 337
rect 778 317 780 322
rect 788 320 790 322
rect 823 325 825 327
rect 833 325 835 329
rect 842 326 844 332
rect 871 339 873 341
rect 876 339 879 341
rect 887 335 889 337
rect 823 317 825 322
rect 833 320 835 322
rect 868 325 870 327
rect 878 325 880 329
rect 887 326 889 332
rect 868 317 870 322
rect 878 320 880 322
rect 16 294 18 296
rect 21 294 24 296
rect 32 290 34 292
rect 13 280 15 282
rect 23 280 25 284
rect 32 281 34 287
rect 61 294 63 296
rect 66 294 69 296
rect 77 290 79 292
rect 13 272 15 277
rect 23 275 25 277
rect 58 280 60 282
rect 68 280 70 284
rect 77 281 79 287
rect 106 294 108 296
rect 111 294 114 296
rect 122 290 124 292
rect 58 272 60 277
rect 68 275 70 277
rect 103 280 105 282
rect 113 280 115 284
rect 122 281 124 287
rect 151 294 153 296
rect 156 294 159 296
rect 167 290 169 292
rect 103 272 105 277
rect 113 275 115 277
rect 148 280 150 282
rect 158 280 160 284
rect 167 281 169 287
rect 196 294 198 296
rect 201 294 204 296
rect 212 290 214 292
rect 148 272 150 277
rect 158 275 160 277
rect 193 280 195 282
rect 203 280 205 284
rect 212 281 214 287
rect 241 294 243 296
rect 246 294 249 296
rect 257 290 259 292
rect 193 272 195 277
rect 203 275 205 277
rect 238 280 240 282
rect 248 280 250 284
rect 257 281 259 287
rect 286 294 288 296
rect 291 294 294 296
rect 302 290 304 292
rect 238 272 240 277
rect 248 275 250 277
rect 283 280 285 282
rect 293 280 295 284
rect 302 281 304 287
rect 331 294 333 296
rect 336 294 339 296
rect 347 290 349 292
rect 283 272 285 277
rect 293 275 295 277
rect 328 280 330 282
rect 338 280 340 284
rect 347 281 349 287
rect 376 294 378 296
rect 381 294 384 296
rect 392 290 394 292
rect 328 272 330 277
rect 338 275 340 277
rect 373 280 375 282
rect 383 280 385 284
rect 392 281 394 287
rect 421 294 423 296
rect 426 294 429 296
rect 437 290 439 292
rect 373 272 375 277
rect 383 275 385 277
rect 418 280 420 282
rect 428 280 430 284
rect 437 281 439 287
rect 466 294 468 296
rect 471 294 474 296
rect 482 290 484 292
rect 418 272 420 277
rect 428 275 430 277
rect 463 280 465 282
rect 473 280 475 284
rect 482 281 484 287
rect 511 294 513 296
rect 516 294 519 296
rect 527 290 529 292
rect 463 272 465 277
rect 473 275 475 277
rect 508 280 510 282
rect 518 280 520 284
rect 527 281 529 287
rect 556 294 558 296
rect 561 294 564 296
rect 572 290 574 292
rect 508 272 510 277
rect 518 275 520 277
rect 553 280 555 282
rect 563 280 565 284
rect 572 281 574 287
rect 601 294 603 296
rect 606 294 609 296
rect 617 290 619 292
rect 553 272 555 277
rect 563 275 565 277
rect 598 280 600 282
rect 608 280 610 284
rect 617 281 619 287
rect 646 294 648 296
rect 651 294 654 296
rect 662 290 664 292
rect 598 272 600 277
rect 608 275 610 277
rect 643 280 645 282
rect 653 280 655 284
rect 662 281 664 287
rect 691 294 693 296
rect 696 294 699 296
rect 707 290 709 292
rect 643 272 645 277
rect 653 275 655 277
rect 688 280 690 282
rect 698 280 700 284
rect 707 281 709 287
rect 736 294 738 296
rect 741 294 744 296
rect 752 290 754 292
rect 688 272 690 277
rect 698 275 700 277
rect 733 280 735 282
rect 743 280 745 284
rect 752 281 754 287
rect 781 294 783 296
rect 786 294 789 296
rect 797 290 799 292
rect 733 272 735 277
rect 743 275 745 277
rect 778 280 780 282
rect 788 280 790 284
rect 797 281 799 287
rect 826 294 828 296
rect 831 294 834 296
rect 842 290 844 292
rect 778 272 780 277
rect 788 275 790 277
rect 823 280 825 282
rect 833 280 835 284
rect 842 281 844 287
rect 871 294 873 296
rect 876 294 879 296
rect 887 290 889 292
rect 823 272 825 277
rect 833 275 835 277
rect 868 280 870 282
rect 878 280 880 284
rect 887 281 889 287
rect 868 272 870 277
rect 878 275 880 277
rect 16 249 18 251
rect 21 249 24 251
rect 32 245 34 247
rect 13 235 15 237
rect 23 235 25 239
rect 32 236 34 242
rect 61 249 63 251
rect 66 249 69 251
rect 77 245 79 247
rect 13 227 15 232
rect 23 230 25 232
rect 58 235 60 237
rect 68 235 70 239
rect 77 236 79 242
rect 106 249 108 251
rect 111 249 114 251
rect 122 245 124 247
rect 58 227 60 232
rect 68 230 70 232
rect 103 235 105 237
rect 113 235 115 239
rect 122 236 124 242
rect 151 249 153 251
rect 156 249 159 251
rect 167 245 169 247
rect 103 227 105 232
rect 113 230 115 232
rect 148 235 150 237
rect 158 235 160 239
rect 167 236 169 242
rect 196 249 198 251
rect 201 249 204 251
rect 212 245 214 247
rect 148 227 150 232
rect 158 230 160 232
rect 193 235 195 237
rect 203 235 205 239
rect 212 236 214 242
rect 241 249 243 251
rect 246 249 249 251
rect 257 245 259 247
rect 193 227 195 232
rect 203 230 205 232
rect 238 235 240 237
rect 248 235 250 239
rect 257 236 259 242
rect 286 249 288 251
rect 291 249 294 251
rect 302 245 304 247
rect 238 227 240 232
rect 248 230 250 232
rect 283 235 285 237
rect 293 235 295 239
rect 302 236 304 242
rect 331 249 333 251
rect 336 249 339 251
rect 347 245 349 247
rect 283 227 285 232
rect 293 230 295 232
rect 328 235 330 237
rect 338 235 340 239
rect 347 236 349 242
rect 376 249 378 251
rect 381 249 384 251
rect 392 245 394 247
rect 328 227 330 232
rect 338 230 340 232
rect 373 235 375 237
rect 383 235 385 239
rect 392 236 394 242
rect 421 249 423 251
rect 426 249 429 251
rect 437 245 439 247
rect 373 227 375 232
rect 383 230 385 232
rect 418 235 420 237
rect 428 235 430 239
rect 437 236 439 242
rect 466 249 468 251
rect 471 249 474 251
rect 482 245 484 247
rect 418 227 420 232
rect 428 230 430 232
rect 463 235 465 237
rect 473 235 475 239
rect 482 236 484 242
rect 511 249 513 251
rect 516 249 519 251
rect 527 245 529 247
rect 463 227 465 232
rect 473 230 475 232
rect 508 235 510 237
rect 518 235 520 239
rect 527 236 529 242
rect 556 249 558 251
rect 561 249 564 251
rect 572 245 574 247
rect 508 227 510 232
rect 518 230 520 232
rect 553 235 555 237
rect 563 235 565 239
rect 572 236 574 242
rect 601 249 603 251
rect 606 249 609 251
rect 617 245 619 247
rect 553 227 555 232
rect 563 230 565 232
rect 598 235 600 237
rect 608 235 610 239
rect 617 236 619 242
rect 646 249 648 251
rect 651 249 654 251
rect 662 245 664 247
rect 598 227 600 232
rect 608 230 610 232
rect 643 235 645 237
rect 653 235 655 239
rect 662 236 664 242
rect 691 249 693 251
rect 696 249 699 251
rect 707 245 709 247
rect 643 227 645 232
rect 653 230 655 232
rect 688 235 690 237
rect 698 235 700 239
rect 707 236 709 242
rect 736 249 738 251
rect 741 249 744 251
rect 752 245 754 247
rect 688 227 690 232
rect 698 230 700 232
rect 733 235 735 237
rect 743 235 745 239
rect 752 236 754 242
rect 781 249 783 251
rect 786 249 789 251
rect 797 245 799 247
rect 733 227 735 232
rect 743 230 745 232
rect 778 235 780 237
rect 788 235 790 239
rect 797 236 799 242
rect 826 249 828 251
rect 831 249 834 251
rect 842 245 844 247
rect 778 227 780 232
rect 788 230 790 232
rect 823 235 825 237
rect 833 235 835 239
rect 842 236 844 242
rect 871 249 873 251
rect 876 249 879 251
rect 887 245 889 247
rect 823 227 825 232
rect 833 230 835 232
rect 868 235 870 237
rect 878 235 880 239
rect 887 236 889 242
rect 868 227 870 232
rect 878 230 880 232
rect 16 204 18 206
rect 21 204 24 206
rect 32 200 34 202
rect 13 190 15 192
rect 23 190 25 194
rect 32 191 34 197
rect 61 204 63 206
rect 66 204 69 206
rect 77 200 79 202
rect 13 182 15 187
rect 23 185 25 187
rect 58 190 60 192
rect 68 190 70 194
rect 77 191 79 197
rect 106 204 108 206
rect 111 204 114 206
rect 122 200 124 202
rect 58 182 60 187
rect 68 185 70 187
rect 103 190 105 192
rect 113 190 115 194
rect 122 191 124 197
rect 151 204 153 206
rect 156 204 159 206
rect 167 200 169 202
rect 103 182 105 187
rect 113 185 115 187
rect 148 190 150 192
rect 158 190 160 194
rect 167 191 169 197
rect 196 204 198 206
rect 201 204 204 206
rect 212 200 214 202
rect 148 182 150 187
rect 158 185 160 187
rect 193 190 195 192
rect 203 190 205 194
rect 212 191 214 197
rect 241 204 243 206
rect 246 204 249 206
rect 257 200 259 202
rect 193 182 195 187
rect 203 185 205 187
rect 238 190 240 192
rect 248 190 250 194
rect 257 191 259 197
rect 286 204 288 206
rect 291 204 294 206
rect 302 200 304 202
rect 238 182 240 187
rect 248 185 250 187
rect 283 190 285 192
rect 293 190 295 194
rect 302 191 304 197
rect 331 204 333 206
rect 336 204 339 206
rect 347 200 349 202
rect 283 182 285 187
rect 293 185 295 187
rect 328 190 330 192
rect 338 190 340 194
rect 347 191 349 197
rect 376 204 378 206
rect 381 204 384 206
rect 392 200 394 202
rect 328 182 330 187
rect 338 185 340 187
rect 373 190 375 192
rect 383 190 385 194
rect 392 191 394 197
rect 421 204 423 206
rect 426 204 429 206
rect 437 200 439 202
rect 373 182 375 187
rect 383 185 385 187
rect 418 190 420 192
rect 428 190 430 194
rect 437 191 439 197
rect 466 204 468 206
rect 471 204 474 206
rect 482 200 484 202
rect 418 182 420 187
rect 428 185 430 187
rect 463 190 465 192
rect 473 190 475 194
rect 482 191 484 197
rect 511 204 513 206
rect 516 204 519 206
rect 527 200 529 202
rect 463 182 465 187
rect 473 185 475 187
rect 508 190 510 192
rect 518 190 520 194
rect 527 191 529 197
rect 556 204 558 206
rect 561 204 564 206
rect 572 200 574 202
rect 508 182 510 187
rect 518 185 520 187
rect 553 190 555 192
rect 563 190 565 194
rect 572 191 574 197
rect 601 204 603 206
rect 606 204 609 206
rect 617 200 619 202
rect 553 182 555 187
rect 563 185 565 187
rect 598 190 600 192
rect 608 190 610 194
rect 617 191 619 197
rect 646 204 648 206
rect 651 204 654 206
rect 662 200 664 202
rect 598 182 600 187
rect 608 185 610 187
rect 643 190 645 192
rect 653 190 655 194
rect 662 191 664 197
rect 691 204 693 206
rect 696 204 699 206
rect 707 200 709 202
rect 643 182 645 187
rect 653 185 655 187
rect 688 190 690 192
rect 698 190 700 194
rect 707 191 709 197
rect 736 204 738 206
rect 741 204 744 206
rect 752 200 754 202
rect 688 182 690 187
rect 698 185 700 187
rect 733 190 735 192
rect 743 190 745 194
rect 752 191 754 197
rect 781 204 783 206
rect 786 204 789 206
rect 797 200 799 202
rect 733 182 735 187
rect 743 185 745 187
rect 778 190 780 192
rect 788 190 790 194
rect 797 191 799 197
rect 826 204 828 206
rect 831 204 834 206
rect 842 200 844 202
rect 778 182 780 187
rect 788 185 790 187
rect 823 190 825 192
rect 833 190 835 194
rect 842 191 844 197
rect 871 204 873 206
rect 876 204 879 206
rect 887 200 889 202
rect 823 182 825 187
rect 833 185 835 187
rect 868 190 870 192
rect 878 190 880 194
rect 887 191 889 197
rect 868 182 870 187
rect 878 185 880 187
rect 16 159 18 161
rect 21 159 24 161
rect 32 155 34 157
rect 13 145 15 147
rect 23 145 25 149
rect 32 146 34 152
rect 61 159 63 161
rect 66 159 69 161
rect 77 155 79 157
rect 13 137 15 142
rect 23 140 25 142
rect 58 145 60 147
rect 68 145 70 149
rect 77 146 79 152
rect 106 159 108 161
rect 111 159 114 161
rect 122 155 124 157
rect 58 137 60 142
rect 68 140 70 142
rect 103 145 105 147
rect 113 145 115 149
rect 122 146 124 152
rect 151 159 153 161
rect 156 159 159 161
rect 167 155 169 157
rect 103 137 105 142
rect 113 140 115 142
rect 148 145 150 147
rect 158 145 160 149
rect 167 146 169 152
rect 196 159 198 161
rect 201 159 204 161
rect 212 155 214 157
rect 148 137 150 142
rect 158 140 160 142
rect 193 145 195 147
rect 203 145 205 149
rect 212 146 214 152
rect 241 159 243 161
rect 246 159 249 161
rect 257 155 259 157
rect 193 137 195 142
rect 203 140 205 142
rect 238 145 240 147
rect 248 145 250 149
rect 257 146 259 152
rect 286 159 288 161
rect 291 159 294 161
rect 302 155 304 157
rect 238 137 240 142
rect 248 140 250 142
rect 283 145 285 147
rect 293 145 295 149
rect 302 146 304 152
rect 331 159 333 161
rect 336 159 339 161
rect 347 155 349 157
rect 283 137 285 142
rect 293 140 295 142
rect 328 145 330 147
rect 338 145 340 149
rect 347 146 349 152
rect 376 159 378 161
rect 381 159 384 161
rect 392 155 394 157
rect 328 137 330 142
rect 338 140 340 142
rect 373 145 375 147
rect 383 145 385 149
rect 392 146 394 152
rect 421 159 423 161
rect 426 159 429 161
rect 437 155 439 157
rect 373 137 375 142
rect 383 140 385 142
rect 418 145 420 147
rect 428 145 430 149
rect 437 146 439 152
rect 466 159 468 161
rect 471 159 474 161
rect 482 155 484 157
rect 418 137 420 142
rect 428 140 430 142
rect 463 145 465 147
rect 473 145 475 149
rect 482 146 484 152
rect 511 159 513 161
rect 516 159 519 161
rect 527 155 529 157
rect 463 137 465 142
rect 473 140 475 142
rect 508 145 510 147
rect 518 145 520 149
rect 527 146 529 152
rect 556 159 558 161
rect 561 159 564 161
rect 572 155 574 157
rect 508 137 510 142
rect 518 140 520 142
rect 553 145 555 147
rect 563 145 565 149
rect 572 146 574 152
rect 601 159 603 161
rect 606 159 609 161
rect 617 155 619 157
rect 553 137 555 142
rect 563 140 565 142
rect 598 145 600 147
rect 608 145 610 149
rect 617 146 619 152
rect 646 159 648 161
rect 651 159 654 161
rect 662 155 664 157
rect 598 137 600 142
rect 608 140 610 142
rect 643 145 645 147
rect 653 145 655 149
rect 662 146 664 152
rect 691 159 693 161
rect 696 159 699 161
rect 707 155 709 157
rect 643 137 645 142
rect 653 140 655 142
rect 688 145 690 147
rect 698 145 700 149
rect 707 146 709 152
rect 736 159 738 161
rect 741 159 744 161
rect 752 155 754 157
rect 688 137 690 142
rect 698 140 700 142
rect 733 145 735 147
rect 743 145 745 149
rect 752 146 754 152
rect 781 159 783 161
rect 786 159 789 161
rect 797 155 799 157
rect 733 137 735 142
rect 743 140 745 142
rect 778 145 780 147
rect 788 145 790 149
rect 797 146 799 152
rect 826 159 828 161
rect 831 159 834 161
rect 842 155 844 157
rect 778 137 780 142
rect 788 140 790 142
rect 823 145 825 147
rect 833 145 835 149
rect 842 146 844 152
rect 871 159 873 161
rect 876 159 879 161
rect 887 155 889 157
rect 823 137 825 142
rect 833 140 835 142
rect 868 145 870 147
rect 878 145 880 149
rect 887 146 889 152
rect 868 137 870 142
rect 878 140 880 142
rect 16 114 18 116
rect 21 114 24 116
rect 32 110 34 112
rect 13 100 15 102
rect 23 100 25 104
rect 32 101 34 107
rect 61 114 63 116
rect 66 114 69 116
rect 77 110 79 112
rect 13 92 15 97
rect 23 95 25 97
rect 58 100 60 102
rect 68 100 70 104
rect 77 101 79 107
rect 106 114 108 116
rect 111 114 114 116
rect 122 110 124 112
rect 58 92 60 97
rect 68 95 70 97
rect 103 100 105 102
rect 113 100 115 104
rect 122 101 124 107
rect 151 114 153 116
rect 156 114 159 116
rect 167 110 169 112
rect 103 92 105 97
rect 113 95 115 97
rect 148 100 150 102
rect 158 100 160 104
rect 167 101 169 107
rect 196 114 198 116
rect 201 114 204 116
rect 212 110 214 112
rect 148 92 150 97
rect 158 95 160 97
rect 193 100 195 102
rect 203 100 205 104
rect 212 101 214 107
rect 241 114 243 116
rect 246 114 249 116
rect 257 110 259 112
rect 193 92 195 97
rect 203 95 205 97
rect 238 100 240 102
rect 248 100 250 104
rect 257 101 259 107
rect 286 114 288 116
rect 291 114 294 116
rect 302 110 304 112
rect 238 92 240 97
rect 248 95 250 97
rect 283 100 285 102
rect 293 100 295 104
rect 302 101 304 107
rect 331 114 333 116
rect 336 114 339 116
rect 347 110 349 112
rect 283 92 285 97
rect 293 95 295 97
rect 328 100 330 102
rect 338 100 340 104
rect 347 101 349 107
rect 376 114 378 116
rect 381 114 384 116
rect 392 110 394 112
rect 328 92 330 97
rect 338 95 340 97
rect 373 100 375 102
rect 383 100 385 104
rect 392 101 394 107
rect 421 114 423 116
rect 426 114 429 116
rect 437 110 439 112
rect 373 92 375 97
rect 383 95 385 97
rect 418 100 420 102
rect 428 100 430 104
rect 437 101 439 107
rect 466 114 468 116
rect 471 114 474 116
rect 482 110 484 112
rect 418 92 420 97
rect 428 95 430 97
rect 463 100 465 102
rect 473 100 475 104
rect 482 101 484 107
rect 511 114 513 116
rect 516 114 519 116
rect 527 110 529 112
rect 463 92 465 97
rect 473 95 475 97
rect 508 100 510 102
rect 518 100 520 104
rect 527 101 529 107
rect 556 114 558 116
rect 561 114 564 116
rect 572 110 574 112
rect 508 92 510 97
rect 518 95 520 97
rect 553 100 555 102
rect 563 100 565 104
rect 572 101 574 107
rect 601 114 603 116
rect 606 114 609 116
rect 617 110 619 112
rect 553 92 555 97
rect 563 95 565 97
rect 598 100 600 102
rect 608 100 610 104
rect 617 101 619 107
rect 646 114 648 116
rect 651 114 654 116
rect 662 110 664 112
rect 598 92 600 97
rect 608 95 610 97
rect 643 100 645 102
rect 653 100 655 104
rect 662 101 664 107
rect 691 114 693 116
rect 696 114 699 116
rect 707 110 709 112
rect 643 92 645 97
rect 653 95 655 97
rect 688 100 690 102
rect 698 100 700 104
rect 707 101 709 107
rect 736 114 738 116
rect 741 114 744 116
rect 752 110 754 112
rect 688 92 690 97
rect 698 95 700 97
rect 733 100 735 102
rect 743 100 745 104
rect 752 101 754 107
rect 781 114 783 116
rect 786 114 789 116
rect 797 110 799 112
rect 733 92 735 97
rect 743 95 745 97
rect 778 100 780 102
rect 788 100 790 104
rect 797 101 799 107
rect 826 114 828 116
rect 831 114 834 116
rect 842 110 844 112
rect 778 92 780 97
rect 788 95 790 97
rect 823 100 825 102
rect 833 100 835 104
rect 842 101 844 107
rect 871 114 873 116
rect 876 114 879 116
rect 887 110 889 112
rect 823 92 825 97
rect 833 95 835 97
rect 868 100 870 102
rect 878 100 880 104
rect 887 101 889 107
rect 868 92 870 97
rect 878 95 880 97
rect 16 69 18 71
rect 21 69 24 71
rect 32 65 34 67
rect 13 55 15 57
rect 23 55 25 59
rect 32 56 34 62
rect 61 69 63 71
rect 66 69 69 71
rect 77 65 79 67
rect 13 47 15 52
rect 23 50 25 52
rect 58 55 60 57
rect 68 55 70 59
rect 77 56 79 62
rect 106 69 108 71
rect 111 69 114 71
rect 122 65 124 67
rect 58 47 60 52
rect 68 50 70 52
rect 103 55 105 57
rect 113 55 115 59
rect 122 56 124 62
rect 151 69 153 71
rect 156 69 159 71
rect 167 65 169 67
rect 103 47 105 52
rect 113 50 115 52
rect 148 55 150 57
rect 158 55 160 59
rect 167 56 169 62
rect 196 69 198 71
rect 201 69 204 71
rect 212 65 214 67
rect 148 47 150 52
rect 158 50 160 52
rect 193 55 195 57
rect 203 55 205 59
rect 212 56 214 62
rect 241 69 243 71
rect 246 69 249 71
rect 257 65 259 67
rect 193 47 195 52
rect 203 50 205 52
rect 238 55 240 57
rect 248 55 250 59
rect 257 56 259 62
rect 286 69 288 71
rect 291 69 294 71
rect 302 65 304 67
rect 238 47 240 52
rect 248 50 250 52
rect 283 55 285 57
rect 293 55 295 59
rect 302 56 304 62
rect 331 69 333 71
rect 336 69 339 71
rect 347 65 349 67
rect 283 47 285 52
rect 293 50 295 52
rect 328 55 330 57
rect 338 55 340 59
rect 347 56 349 62
rect 376 69 378 71
rect 381 69 384 71
rect 392 65 394 67
rect 328 47 330 52
rect 338 50 340 52
rect 373 55 375 57
rect 383 55 385 59
rect 392 56 394 62
rect 421 69 423 71
rect 426 69 429 71
rect 437 65 439 67
rect 373 47 375 52
rect 383 50 385 52
rect 418 55 420 57
rect 428 55 430 59
rect 437 56 439 62
rect 466 69 468 71
rect 471 69 474 71
rect 482 65 484 67
rect 418 47 420 52
rect 428 50 430 52
rect 463 55 465 57
rect 473 55 475 59
rect 482 56 484 62
rect 511 69 513 71
rect 516 69 519 71
rect 527 65 529 67
rect 463 47 465 52
rect 473 50 475 52
rect 508 55 510 57
rect 518 55 520 59
rect 527 56 529 62
rect 556 69 558 71
rect 561 69 564 71
rect 572 65 574 67
rect 508 47 510 52
rect 518 50 520 52
rect 553 55 555 57
rect 563 55 565 59
rect 572 56 574 62
rect 601 69 603 71
rect 606 69 609 71
rect 617 65 619 67
rect 553 47 555 52
rect 563 50 565 52
rect 598 55 600 57
rect 608 55 610 59
rect 617 56 619 62
rect 646 69 648 71
rect 651 69 654 71
rect 662 65 664 67
rect 598 47 600 52
rect 608 50 610 52
rect 643 55 645 57
rect 653 55 655 59
rect 662 56 664 62
rect 691 69 693 71
rect 696 69 699 71
rect 707 65 709 67
rect 643 47 645 52
rect 653 50 655 52
rect 688 55 690 57
rect 698 55 700 59
rect 707 56 709 62
rect 736 69 738 71
rect 741 69 744 71
rect 752 65 754 67
rect 688 47 690 52
rect 698 50 700 52
rect 733 55 735 57
rect 743 55 745 59
rect 752 56 754 62
rect 781 69 783 71
rect 786 69 789 71
rect 797 65 799 67
rect 733 47 735 52
rect 743 50 745 52
rect 778 55 780 57
rect 788 55 790 59
rect 797 56 799 62
rect 826 69 828 71
rect 831 69 834 71
rect 842 65 844 67
rect 778 47 780 52
rect 788 50 790 52
rect 823 55 825 57
rect 833 55 835 59
rect 842 56 844 62
rect 871 69 873 71
rect 876 69 879 71
rect 887 65 889 67
rect 823 47 825 52
rect 833 50 835 52
rect 868 55 870 57
rect 878 55 880 59
rect 887 56 889 62
rect 868 47 870 52
rect 878 50 880 52
rect 16 24 18 26
rect 21 24 24 26
rect 32 20 34 22
rect 13 10 15 12
rect 23 10 25 14
rect 32 11 34 17
rect 61 24 63 26
rect 66 24 69 26
rect 77 20 79 22
rect 13 2 15 7
rect 23 5 25 7
rect 58 10 60 12
rect 68 10 70 14
rect 77 11 79 17
rect 106 24 108 26
rect 111 24 114 26
rect 122 20 124 22
rect 58 2 60 7
rect 68 5 70 7
rect 103 10 105 12
rect 113 10 115 14
rect 122 11 124 17
rect 151 24 153 26
rect 156 24 159 26
rect 167 20 169 22
rect 103 2 105 7
rect 113 5 115 7
rect 148 10 150 12
rect 158 10 160 14
rect 167 11 169 17
rect 196 24 198 26
rect 201 24 204 26
rect 212 20 214 22
rect 148 2 150 7
rect 158 5 160 7
rect 193 10 195 12
rect 203 10 205 14
rect 212 11 214 17
rect 241 24 243 26
rect 246 24 249 26
rect 257 20 259 22
rect 193 2 195 7
rect 203 5 205 7
rect 238 10 240 12
rect 248 10 250 14
rect 257 11 259 17
rect 286 24 288 26
rect 291 24 294 26
rect 302 20 304 22
rect 238 2 240 7
rect 248 5 250 7
rect 283 10 285 12
rect 293 10 295 14
rect 302 11 304 17
rect 331 24 333 26
rect 336 24 339 26
rect 347 20 349 22
rect 283 2 285 7
rect 293 5 295 7
rect 328 10 330 12
rect 338 10 340 14
rect 347 11 349 17
rect 376 24 378 26
rect 381 24 384 26
rect 392 20 394 22
rect 328 2 330 7
rect 338 5 340 7
rect 373 10 375 12
rect 383 10 385 14
rect 392 11 394 17
rect 421 24 423 26
rect 426 24 429 26
rect 437 20 439 22
rect 373 2 375 7
rect 383 5 385 7
rect 418 10 420 12
rect 428 10 430 14
rect 437 11 439 17
rect 466 24 468 26
rect 471 24 474 26
rect 482 20 484 22
rect 418 2 420 7
rect 428 5 430 7
rect 463 10 465 12
rect 473 10 475 14
rect 482 11 484 17
rect 511 24 513 26
rect 516 24 519 26
rect 527 20 529 22
rect 463 2 465 7
rect 473 5 475 7
rect 508 10 510 12
rect 518 10 520 14
rect 527 11 529 17
rect 556 24 558 26
rect 561 24 564 26
rect 572 20 574 22
rect 508 2 510 7
rect 518 5 520 7
rect 553 10 555 12
rect 563 10 565 14
rect 572 11 574 17
rect 601 24 603 26
rect 606 24 609 26
rect 617 20 619 22
rect 553 2 555 7
rect 563 5 565 7
rect 598 10 600 12
rect 608 10 610 14
rect 617 11 619 17
rect 646 24 648 26
rect 651 24 654 26
rect 662 20 664 22
rect 598 2 600 7
rect 608 5 610 7
rect 643 10 645 12
rect 653 10 655 14
rect 662 11 664 17
rect 691 24 693 26
rect 696 24 699 26
rect 707 20 709 22
rect 643 2 645 7
rect 653 5 655 7
rect 688 10 690 12
rect 698 10 700 14
rect 707 11 709 17
rect 736 24 738 26
rect 741 24 744 26
rect 752 20 754 22
rect 688 2 690 7
rect 698 5 700 7
rect 733 10 735 12
rect 743 10 745 14
rect 752 11 754 17
rect 781 24 783 26
rect 786 24 789 26
rect 797 20 799 22
rect 733 2 735 7
rect 743 5 745 7
rect 778 10 780 12
rect 788 10 790 14
rect 797 11 799 17
rect 826 24 828 26
rect 831 24 834 26
rect 842 20 844 22
rect 778 2 780 7
rect 788 5 790 7
rect 823 10 825 12
rect 833 10 835 14
rect 842 11 844 17
rect 871 24 873 26
rect 876 24 879 26
rect 887 20 889 22
rect 823 2 825 7
rect 833 5 835 7
rect 868 10 870 12
rect 878 10 880 14
rect 887 11 889 17
rect 868 2 870 7
rect 878 5 880 7
rect -292 -163 -290 -159
rect -287 -163 -285 -161
rect -271 -165 -268 -163
rect -263 -165 -261 -163
rect -292 -171 -290 -169
rect -287 -171 -285 -169
rect -200 -157 -198 -155
rect -195 -157 -192 -155
rect -184 -161 -182 -159
rect -260 -170 -258 -168
rect -287 -175 -286 -171
rect -203 -171 -201 -169
rect -193 -171 -191 -167
rect -184 -170 -182 -164
rect -260 -178 -258 -176
rect -203 -179 -201 -174
rect -193 -176 -191 -174
<< polycontact >>
rect 24 878 28 882
rect 19 867 23 871
rect 69 878 73 882
rect 34 865 38 869
rect 64 867 68 871
rect 15 856 19 860
rect 114 878 118 882
rect 79 865 83 869
rect 109 867 113 871
rect 60 856 64 860
rect 159 878 163 882
rect 124 865 128 869
rect 154 867 158 871
rect 105 856 109 860
rect 204 878 208 882
rect 169 865 173 869
rect 199 867 203 871
rect 150 856 154 860
rect 249 878 253 882
rect 214 865 218 869
rect 244 867 248 871
rect 195 856 199 860
rect 294 878 298 882
rect 259 865 263 869
rect 289 867 293 871
rect 240 856 244 860
rect 339 878 343 882
rect 304 865 308 869
rect 334 867 338 871
rect 285 856 289 860
rect 384 878 388 882
rect 349 865 353 869
rect 379 867 383 871
rect 330 856 334 860
rect 429 878 433 882
rect 394 865 398 869
rect 424 867 428 871
rect 375 856 379 860
rect 474 878 478 882
rect 439 865 443 869
rect 469 867 473 871
rect 420 856 424 860
rect 519 878 523 882
rect 484 865 488 869
rect 514 867 518 871
rect 465 856 469 860
rect 564 878 568 882
rect 529 865 533 869
rect 559 867 563 871
rect 510 856 514 860
rect 609 878 613 882
rect 574 865 578 869
rect 604 867 608 871
rect 555 856 559 860
rect 654 878 658 882
rect 619 865 623 869
rect 649 867 653 871
rect 600 856 604 860
rect 699 878 703 882
rect 664 865 668 869
rect 694 867 698 871
rect 645 856 649 860
rect 744 878 748 882
rect 709 865 713 869
rect 739 867 743 871
rect 690 856 694 860
rect 789 878 793 882
rect 754 865 758 869
rect 784 867 788 871
rect 735 856 739 860
rect 834 878 838 882
rect 799 865 803 869
rect 829 867 833 871
rect 780 856 784 860
rect 879 878 883 882
rect 844 865 848 869
rect 874 867 878 871
rect 825 856 829 860
rect 889 865 893 869
rect 870 856 874 860
rect 24 833 28 837
rect 19 822 23 826
rect 69 833 73 837
rect 34 820 38 824
rect 64 822 68 826
rect 15 811 19 815
rect 114 833 118 837
rect 79 820 83 824
rect 109 822 113 826
rect 60 811 64 815
rect 159 833 163 837
rect 124 820 128 824
rect 154 822 158 826
rect 105 811 109 815
rect 204 833 208 837
rect 169 820 173 824
rect 199 822 203 826
rect 150 811 154 815
rect 249 833 253 837
rect 214 820 218 824
rect 244 822 248 826
rect 195 811 199 815
rect 294 833 298 837
rect 259 820 263 824
rect 289 822 293 826
rect 240 811 244 815
rect 339 833 343 837
rect 304 820 308 824
rect 334 822 338 826
rect 285 811 289 815
rect 384 833 388 837
rect 349 820 353 824
rect 379 822 383 826
rect 330 811 334 815
rect 429 833 433 837
rect 394 820 398 824
rect 424 822 428 826
rect 375 811 379 815
rect 474 833 478 837
rect 439 820 443 824
rect 469 822 473 826
rect 420 811 424 815
rect 519 833 523 837
rect 484 820 488 824
rect 514 822 518 826
rect 465 811 469 815
rect 564 833 568 837
rect 529 820 533 824
rect 559 822 563 826
rect 510 811 514 815
rect 609 833 613 837
rect 574 820 578 824
rect 604 822 608 826
rect 555 811 559 815
rect 654 833 658 837
rect 619 820 623 824
rect 649 822 653 826
rect 600 811 604 815
rect 699 833 703 837
rect 664 820 668 824
rect 694 822 698 826
rect 645 811 649 815
rect 744 833 748 837
rect 709 820 713 824
rect 739 822 743 826
rect 690 811 694 815
rect 789 833 793 837
rect 754 820 758 824
rect 784 822 788 826
rect 735 811 739 815
rect 834 833 838 837
rect 799 820 803 824
rect 829 822 833 826
rect 780 811 784 815
rect 879 833 883 837
rect 844 820 848 824
rect 874 822 878 826
rect 825 811 829 815
rect 889 820 893 824
rect 870 811 874 815
rect 24 788 28 792
rect 19 777 23 781
rect 69 788 73 792
rect 34 775 38 779
rect 64 777 68 781
rect 15 766 19 770
rect 114 788 118 792
rect 79 775 83 779
rect 109 777 113 781
rect 60 766 64 770
rect 159 788 163 792
rect 124 775 128 779
rect 154 777 158 781
rect 105 766 109 770
rect 204 788 208 792
rect 169 775 173 779
rect 199 777 203 781
rect 150 766 154 770
rect 249 788 253 792
rect 214 775 218 779
rect 244 777 248 781
rect 195 766 199 770
rect 294 788 298 792
rect 259 775 263 779
rect 289 777 293 781
rect 240 766 244 770
rect 339 788 343 792
rect 304 775 308 779
rect 334 777 338 781
rect 285 766 289 770
rect 384 788 388 792
rect 349 775 353 779
rect 379 777 383 781
rect 330 766 334 770
rect 429 788 433 792
rect 394 775 398 779
rect 424 777 428 781
rect 375 766 379 770
rect 474 788 478 792
rect 439 775 443 779
rect 469 777 473 781
rect 420 766 424 770
rect 519 788 523 792
rect 484 775 488 779
rect 514 777 518 781
rect 465 766 469 770
rect 564 788 568 792
rect 529 775 533 779
rect 559 777 563 781
rect 510 766 514 770
rect 609 788 613 792
rect 574 775 578 779
rect 604 777 608 781
rect 555 766 559 770
rect 654 788 658 792
rect 619 775 623 779
rect 649 777 653 781
rect 600 766 604 770
rect 699 788 703 792
rect 664 775 668 779
rect 694 777 698 781
rect 645 766 649 770
rect 744 788 748 792
rect 709 775 713 779
rect 739 777 743 781
rect 690 766 694 770
rect 789 788 793 792
rect 754 775 758 779
rect 784 777 788 781
rect 735 766 739 770
rect 834 788 838 792
rect 799 775 803 779
rect 829 777 833 781
rect 780 766 784 770
rect 879 788 883 792
rect 844 775 848 779
rect 874 777 878 781
rect 825 766 829 770
rect 889 775 893 779
rect 870 766 874 770
rect 24 743 28 747
rect 19 732 23 736
rect 69 743 73 747
rect 34 730 38 734
rect 64 732 68 736
rect 15 721 19 725
rect 114 743 118 747
rect 79 730 83 734
rect 109 732 113 736
rect 60 721 64 725
rect 159 743 163 747
rect 124 730 128 734
rect 154 732 158 736
rect 105 721 109 725
rect 204 743 208 747
rect 169 730 173 734
rect 199 732 203 736
rect 150 721 154 725
rect 249 743 253 747
rect 214 730 218 734
rect 244 732 248 736
rect 195 721 199 725
rect 294 743 298 747
rect 259 730 263 734
rect 289 732 293 736
rect 240 721 244 725
rect 339 743 343 747
rect 304 730 308 734
rect 334 732 338 736
rect 285 721 289 725
rect 384 743 388 747
rect 349 730 353 734
rect 379 732 383 736
rect 330 721 334 725
rect 429 743 433 747
rect 394 730 398 734
rect 424 732 428 736
rect 375 721 379 725
rect 474 743 478 747
rect 439 730 443 734
rect 469 732 473 736
rect 420 721 424 725
rect 519 743 523 747
rect 484 730 488 734
rect 514 732 518 736
rect 465 721 469 725
rect 564 743 568 747
rect 529 730 533 734
rect 559 732 563 736
rect 510 721 514 725
rect 609 743 613 747
rect 574 730 578 734
rect 604 732 608 736
rect 555 721 559 725
rect 654 743 658 747
rect 619 730 623 734
rect 649 732 653 736
rect 600 721 604 725
rect 699 743 703 747
rect 664 730 668 734
rect 694 732 698 736
rect 645 721 649 725
rect 744 743 748 747
rect 709 730 713 734
rect 739 732 743 736
rect 690 721 694 725
rect 789 743 793 747
rect 754 730 758 734
rect 784 732 788 736
rect 735 721 739 725
rect 834 743 838 747
rect 799 730 803 734
rect 829 732 833 736
rect 780 721 784 725
rect 879 743 883 747
rect 844 730 848 734
rect 874 732 878 736
rect 825 721 829 725
rect 889 730 893 734
rect 870 721 874 725
rect 24 698 28 702
rect 19 687 23 691
rect 69 698 73 702
rect 34 685 38 689
rect 64 687 68 691
rect 15 676 19 680
rect 114 698 118 702
rect 79 685 83 689
rect 109 687 113 691
rect 60 676 64 680
rect 159 698 163 702
rect 124 685 128 689
rect 154 687 158 691
rect 105 676 109 680
rect 204 698 208 702
rect 169 685 173 689
rect 199 687 203 691
rect 150 676 154 680
rect 249 698 253 702
rect 214 685 218 689
rect 244 687 248 691
rect 195 676 199 680
rect 294 698 298 702
rect 259 685 263 689
rect 289 687 293 691
rect 240 676 244 680
rect 339 698 343 702
rect 304 685 308 689
rect 334 687 338 691
rect 285 676 289 680
rect 384 698 388 702
rect 349 685 353 689
rect 379 687 383 691
rect 330 676 334 680
rect 429 698 433 702
rect 394 685 398 689
rect 424 687 428 691
rect 375 676 379 680
rect 474 698 478 702
rect 439 685 443 689
rect 469 687 473 691
rect 420 676 424 680
rect 519 698 523 702
rect 484 685 488 689
rect 514 687 518 691
rect 465 676 469 680
rect 564 698 568 702
rect 529 685 533 689
rect 559 687 563 691
rect 510 676 514 680
rect 609 698 613 702
rect 574 685 578 689
rect 604 687 608 691
rect 555 676 559 680
rect 654 698 658 702
rect 619 685 623 689
rect 649 687 653 691
rect 600 676 604 680
rect 699 698 703 702
rect 664 685 668 689
rect 694 687 698 691
rect 645 676 649 680
rect 744 698 748 702
rect 709 685 713 689
rect 739 687 743 691
rect 690 676 694 680
rect 789 698 793 702
rect 754 685 758 689
rect 784 687 788 691
rect 735 676 739 680
rect 834 698 838 702
rect 799 685 803 689
rect 829 687 833 691
rect 780 676 784 680
rect 879 698 883 702
rect 844 685 848 689
rect 874 687 878 691
rect 825 676 829 680
rect 889 685 893 689
rect 870 676 874 680
rect 24 653 28 657
rect 19 642 23 646
rect 69 653 73 657
rect 34 640 38 644
rect 64 642 68 646
rect 15 631 19 635
rect 114 653 118 657
rect 79 640 83 644
rect 109 642 113 646
rect 60 631 64 635
rect 159 653 163 657
rect 124 640 128 644
rect 154 642 158 646
rect 105 631 109 635
rect 204 653 208 657
rect 169 640 173 644
rect 199 642 203 646
rect 150 631 154 635
rect 249 653 253 657
rect 214 640 218 644
rect 244 642 248 646
rect 195 631 199 635
rect 294 653 298 657
rect 259 640 263 644
rect 289 642 293 646
rect 240 631 244 635
rect 339 653 343 657
rect 304 640 308 644
rect 334 642 338 646
rect 285 631 289 635
rect 384 653 388 657
rect 349 640 353 644
rect 379 642 383 646
rect 330 631 334 635
rect 429 653 433 657
rect 394 640 398 644
rect 424 642 428 646
rect 375 631 379 635
rect 474 653 478 657
rect 439 640 443 644
rect 469 642 473 646
rect 420 631 424 635
rect 519 653 523 657
rect 484 640 488 644
rect 514 642 518 646
rect 465 631 469 635
rect 564 653 568 657
rect 529 640 533 644
rect 559 642 563 646
rect 510 631 514 635
rect 609 653 613 657
rect 574 640 578 644
rect 604 642 608 646
rect 555 631 559 635
rect 654 653 658 657
rect 619 640 623 644
rect 649 642 653 646
rect 600 631 604 635
rect 699 653 703 657
rect 664 640 668 644
rect 694 642 698 646
rect 645 631 649 635
rect 744 653 748 657
rect 709 640 713 644
rect 739 642 743 646
rect 690 631 694 635
rect 789 653 793 657
rect 754 640 758 644
rect 784 642 788 646
rect 735 631 739 635
rect 834 653 838 657
rect 799 640 803 644
rect 829 642 833 646
rect 780 631 784 635
rect 879 653 883 657
rect 844 640 848 644
rect 874 642 878 646
rect 825 631 829 635
rect 889 640 893 644
rect 870 631 874 635
rect 24 608 28 612
rect 19 597 23 601
rect 69 608 73 612
rect 34 595 38 599
rect 64 597 68 601
rect 15 586 19 590
rect 114 608 118 612
rect 79 595 83 599
rect 109 597 113 601
rect 60 586 64 590
rect 159 608 163 612
rect 124 595 128 599
rect 154 597 158 601
rect 105 586 109 590
rect 204 608 208 612
rect 169 595 173 599
rect 199 597 203 601
rect 150 586 154 590
rect 249 608 253 612
rect 214 595 218 599
rect 244 597 248 601
rect 195 586 199 590
rect 294 608 298 612
rect 259 595 263 599
rect 289 597 293 601
rect 240 586 244 590
rect 339 608 343 612
rect 304 595 308 599
rect 334 597 338 601
rect 285 586 289 590
rect 384 608 388 612
rect 349 595 353 599
rect 379 597 383 601
rect 330 586 334 590
rect 429 608 433 612
rect 394 595 398 599
rect 424 597 428 601
rect 375 586 379 590
rect 474 608 478 612
rect 439 595 443 599
rect 469 597 473 601
rect 420 586 424 590
rect 519 608 523 612
rect 484 595 488 599
rect 514 597 518 601
rect 465 586 469 590
rect 564 608 568 612
rect 529 595 533 599
rect 559 597 563 601
rect 510 586 514 590
rect 609 608 613 612
rect 574 595 578 599
rect 604 597 608 601
rect 555 586 559 590
rect 654 608 658 612
rect 619 595 623 599
rect 649 597 653 601
rect 600 586 604 590
rect 699 608 703 612
rect 664 595 668 599
rect 694 597 698 601
rect 645 586 649 590
rect 744 608 748 612
rect 709 595 713 599
rect 739 597 743 601
rect 690 586 694 590
rect 789 608 793 612
rect 754 595 758 599
rect 784 597 788 601
rect 735 586 739 590
rect 834 608 838 612
rect 799 595 803 599
rect 829 597 833 601
rect 780 586 784 590
rect 879 608 883 612
rect 844 595 848 599
rect 874 597 878 601
rect 825 586 829 590
rect 889 595 893 599
rect 870 586 874 590
rect 24 563 28 567
rect 19 552 23 556
rect 69 563 73 567
rect 34 550 38 554
rect 64 552 68 556
rect 15 541 19 545
rect 114 563 118 567
rect 79 550 83 554
rect 109 552 113 556
rect 60 541 64 545
rect 159 563 163 567
rect 124 550 128 554
rect 154 552 158 556
rect 105 541 109 545
rect 204 563 208 567
rect 169 550 173 554
rect 199 552 203 556
rect 150 541 154 545
rect 249 563 253 567
rect 214 550 218 554
rect 244 552 248 556
rect 195 541 199 545
rect 294 563 298 567
rect 259 550 263 554
rect 289 552 293 556
rect 240 541 244 545
rect 339 563 343 567
rect 304 550 308 554
rect 334 552 338 556
rect 285 541 289 545
rect 384 563 388 567
rect 349 550 353 554
rect 379 552 383 556
rect 330 541 334 545
rect 429 563 433 567
rect 394 550 398 554
rect 424 552 428 556
rect 375 541 379 545
rect 474 563 478 567
rect 439 550 443 554
rect 469 552 473 556
rect 420 541 424 545
rect 519 563 523 567
rect 484 550 488 554
rect 514 552 518 556
rect 465 541 469 545
rect 564 563 568 567
rect 529 550 533 554
rect 559 552 563 556
rect 510 541 514 545
rect 609 563 613 567
rect 574 550 578 554
rect 604 552 608 556
rect 555 541 559 545
rect 654 563 658 567
rect 619 550 623 554
rect 649 552 653 556
rect 600 541 604 545
rect 699 563 703 567
rect 664 550 668 554
rect 694 552 698 556
rect 645 541 649 545
rect 744 563 748 567
rect 709 550 713 554
rect 739 552 743 556
rect 690 541 694 545
rect 789 563 793 567
rect 754 550 758 554
rect 784 552 788 556
rect 735 541 739 545
rect 834 563 838 567
rect 799 550 803 554
rect 829 552 833 556
rect 780 541 784 545
rect 879 563 883 567
rect 844 550 848 554
rect 874 552 878 556
rect 825 541 829 545
rect 889 550 893 554
rect 870 541 874 545
rect 24 518 28 522
rect 19 507 23 511
rect 69 518 73 522
rect 34 505 38 509
rect 64 507 68 511
rect 15 496 19 500
rect 114 518 118 522
rect 79 505 83 509
rect 109 507 113 511
rect 60 496 64 500
rect 159 518 163 522
rect 124 505 128 509
rect 154 507 158 511
rect 105 496 109 500
rect 204 518 208 522
rect 169 505 173 509
rect 199 507 203 511
rect 150 496 154 500
rect 249 518 253 522
rect 214 505 218 509
rect 244 507 248 511
rect 195 496 199 500
rect 294 518 298 522
rect 259 505 263 509
rect 289 507 293 511
rect 240 496 244 500
rect 339 518 343 522
rect 304 505 308 509
rect 334 507 338 511
rect 285 496 289 500
rect 384 518 388 522
rect 349 505 353 509
rect 379 507 383 511
rect 330 496 334 500
rect 429 518 433 522
rect 394 505 398 509
rect 424 507 428 511
rect 375 496 379 500
rect 474 518 478 522
rect 439 505 443 509
rect 469 507 473 511
rect 420 496 424 500
rect 519 518 523 522
rect 484 505 488 509
rect 514 507 518 511
rect 465 496 469 500
rect 564 518 568 522
rect 529 505 533 509
rect 559 507 563 511
rect 510 496 514 500
rect 609 518 613 522
rect 574 505 578 509
rect 604 507 608 511
rect 555 496 559 500
rect 654 518 658 522
rect 619 505 623 509
rect 649 507 653 511
rect 600 496 604 500
rect 699 518 703 522
rect 664 505 668 509
rect 694 507 698 511
rect 645 496 649 500
rect 744 518 748 522
rect 709 505 713 509
rect 739 507 743 511
rect 690 496 694 500
rect 789 518 793 522
rect 754 505 758 509
rect 784 507 788 511
rect 735 496 739 500
rect 834 518 838 522
rect 799 505 803 509
rect 829 507 833 511
rect 780 496 784 500
rect 879 518 883 522
rect 844 505 848 509
rect 874 507 878 511
rect 825 496 829 500
rect 889 505 893 509
rect 870 496 874 500
rect 24 473 28 477
rect 19 462 23 466
rect 69 473 73 477
rect 34 460 38 464
rect 64 462 68 466
rect 15 451 19 455
rect 114 473 118 477
rect 79 460 83 464
rect 109 462 113 466
rect 60 451 64 455
rect 159 473 163 477
rect 124 460 128 464
rect 154 462 158 466
rect 105 451 109 455
rect 204 473 208 477
rect 169 460 173 464
rect 199 462 203 466
rect 150 451 154 455
rect 249 473 253 477
rect 214 460 218 464
rect 244 462 248 466
rect 195 451 199 455
rect 294 473 298 477
rect 259 460 263 464
rect 289 462 293 466
rect 240 451 244 455
rect 339 473 343 477
rect 304 460 308 464
rect 334 462 338 466
rect 285 451 289 455
rect 384 473 388 477
rect 349 460 353 464
rect 379 462 383 466
rect 330 451 334 455
rect 429 473 433 477
rect 394 460 398 464
rect 424 462 428 466
rect 375 451 379 455
rect 474 473 478 477
rect 439 460 443 464
rect 469 462 473 466
rect 420 451 424 455
rect 519 473 523 477
rect 484 460 488 464
rect 514 462 518 466
rect 465 451 469 455
rect 564 473 568 477
rect 529 460 533 464
rect 559 462 563 466
rect 510 451 514 455
rect 609 473 613 477
rect 574 460 578 464
rect 604 462 608 466
rect 555 451 559 455
rect 654 473 658 477
rect 619 460 623 464
rect 649 462 653 466
rect 600 451 604 455
rect 699 473 703 477
rect 664 460 668 464
rect 694 462 698 466
rect 645 451 649 455
rect 744 473 748 477
rect 709 460 713 464
rect 739 462 743 466
rect 690 451 694 455
rect 789 473 793 477
rect 754 460 758 464
rect 784 462 788 466
rect 735 451 739 455
rect 834 473 838 477
rect 799 460 803 464
rect 829 462 833 466
rect 780 451 784 455
rect 879 473 883 477
rect 844 460 848 464
rect 874 462 878 466
rect 825 451 829 455
rect 889 460 893 464
rect 870 451 874 455
rect 24 428 28 432
rect 19 417 23 421
rect 69 428 73 432
rect 34 415 38 419
rect 64 417 68 421
rect 15 406 19 410
rect 114 428 118 432
rect 79 415 83 419
rect 109 417 113 421
rect 60 406 64 410
rect 159 428 163 432
rect 124 415 128 419
rect 154 417 158 421
rect 105 406 109 410
rect 204 428 208 432
rect 169 415 173 419
rect 199 417 203 421
rect 150 406 154 410
rect 249 428 253 432
rect 214 415 218 419
rect 244 417 248 421
rect 195 406 199 410
rect 294 428 298 432
rect 259 415 263 419
rect 289 417 293 421
rect 240 406 244 410
rect 339 428 343 432
rect 304 415 308 419
rect 334 417 338 421
rect 285 406 289 410
rect 384 428 388 432
rect 349 415 353 419
rect 379 417 383 421
rect 330 406 334 410
rect 429 428 433 432
rect 394 415 398 419
rect 424 417 428 421
rect 375 406 379 410
rect 474 428 478 432
rect 439 415 443 419
rect 469 417 473 421
rect 420 406 424 410
rect 519 428 523 432
rect 484 415 488 419
rect 514 417 518 421
rect 465 406 469 410
rect 564 428 568 432
rect 529 415 533 419
rect 559 417 563 421
rect 510 406 514 410
rect 609 428 613 432
rect 574 415 578 419
rect 604 417 608 421
rect 555 406 559 410
rect 654 428 658 432
rect 619 415 623 419
rect 649 417 653 421
rect 600 406 604 410
rect 699 428 703 432
rect 664 415 668 419
rect 694 417 698 421
rect 645 406 649 410
rect 744 428 748 432
rect 709 415 713 419
rect 739 417 743 421
rect 690 406 694 410
rect 789 428 793 432
rect 754 415 758 419
rect 784 417 788 421
rect 735 406 739 410
rect 834 428 838 432
rect 799 415 803 419
rect 829 417 833 421
rect 780 406 784 410
rect 879 428 883 432
rect 844 415 848 419
rect 874 417 878 421
rect 825 406 829 410
rect 889 415 893 419
rect 870 406 874 410
rect 24 383 28 387
rect 19 372 23 376
rect 69 383 73 387
rect 34 370 38 374
rect 64 372 68 376
rect 15 361 19 365
rect 114 383 118 387
rect 79 370 83 374
rect 109 372 113 376
rect 60 361 64 365
rect 159 383 163 387
rect 124 370 128 374
rect 154 372 158 376
rect 105 361 109 365
rect 204 383 208 387
rect 169 370 173 374
rect 199 372 203 376
rect 150 361 154 365
rect 249 383 253 387
rect 214 370 218 374
rect 244 372 248 376
rect 195 361 199 365
rect 294 383 298 387
rect 259 370 263 374
rect 289 372 293 376
rect 240 361 244 365
rect 339 383 343 387
rect 304 370 308 374
rect 334 372 338 376
rect 285 361 289 365
rect 384 383 388 387
rect 349 370 353 374
rect 379 372 383 376
rect 330 361 334 365
rect 429 383 433 387
rect 394 370 398 374
rect 424 372 428 376
rect 375 361 379 365
rect 474 383 478 387
rect 439 370 443 374
rect 469 372 473 376
rect 420 361 424 365
rect 519 383 523 387
rect 484 370 488 374
rect 514 372 518 376
rect 465 361 469 365
rect 564 383 568 387
rect 529 370 533 374
rect 559 372 563 376
rect 510 361 514 365
rect 609 383 613 387
rect 574 370 578 374
rect 604 372 608 376
rect 555 361 559 365
rect 654 383 658 387
rect 619 370 623 374
rect 649 372 653 376
rect 600 361 604 365
rect 699 383 703 387
rect 664 370 668 374
rect 694 372 698 376
rect 645 361 649 365
rect 744 383 748 387
rect 709 370 713 374
rect 739 372 743 376
rect 690 361 694 365
rect 789 383 793 387
rect 754 370 758 374
rect 784 372 788 376
rect 735 361 739 365
rect 834 383 838 387
rect 799 370 803 374
rect 829 372 833 376
rect 780 361 784 365
rect 879 383 883 387
rect 844 370 848 374
rect 874 372 878 376
rect 825 361 829 365
rect 889 370 893 374
rect 870 361 874 365
rect 24 338 28 342
rect 19 327 23 331
rect 69 338 73 342
rect 34 325 38 329
rect 64 327 68 331
rect 15 316 19 320
rect 114 338 118 342
rect 79 325 83 329
rect 109 327 113 331
rect 60 316 64 320
rect 159 338 163 342
rect 124 325 128 329
rect 154 327 158 331
rect 105 316 109 320
rect 204 338 208 342
rect 169 325 173 329
rect 199 327 203 331
rect 150 316 154 320
rect 249 338 253 342
rect 214 325 218 329
rect 244 327 248 331
rect 195 316 199 320
rect 294 338 298 342
rect 259 325 263 329
rect 289 327 293 331
rect 240 316 244 320
rect 339 338 343 342
rect 304 325 308 329
rect 334 327 338 331
rect 285 316 289 320
rect 384 338 388 342
rect 349 325 353 329
rect 379 327 383 331
rect 330 316 334 320
rect 429 338 433 342
rect 394 325 398 329
rect 424 327 428 331
rect 375 316 379 320
rect 474 338 478 342
rect 439 325 443 329
rect 469 327 473 331
rect 420 316 424 320
rect 519 338 523 342
rect 484 325 488 329
rect 514 327 518 331
rect 465 316 469 320
rect 564 338 568 342
rect 529 325 533 329
rect 559 327 563 331
rect 510 316 514 320
rect 609 338 613 342
rect 574 325 578 329
rect 604 327 608 331
rect 555 316 559 320
rect 654 338 658 342
rect 619 325 623 329
rect 649 327 653 331
rect 600 316 604 320
rect 699 338 703 342
rect 664 325 668 329
rect 694 327 698 331
rect 645 316 649 320
rect 744 338 748 342
rect 709 325 713 329
rect 739 327 743 331
rect 690 316 694 320
rect 789 338 793 342
rect 754 325 758 329
rect 784 327 788 331
rect 735 316 739 320
rect 834 338 838 342
rect 799 325 803 329
rect 829 327 833 331
rect 780 316 784 320
rect 879 338 883 342
rect 844 325 848 329
rect 874 327 878 331
rect 825 316 829 320
rect 889 325 893 329
rect 870 316 874 320
rect 24 293 28 297
rect 19 282 23 286
rect 69 293 73 297
rect 34 280 38 284
rect 64 282 68 286
rect 15 271 19 275
rect 114 293 118 297
rect 79 280 83 284
rect 109 282 113 286
rect 60 271 64 275
rect 159 293 163 297
rect 124 280 128 284
rect 154 282 158 286
rect 105 271 109 275
rect 204 293 208 297
rect 169 280 173 284
rect 199 282 203 286
rect 150 271 154 275
rect 249 293 253 297
rect 214 280 218 284
rect 244 282 248 286
rect 195 271 199 275
rect 294 293 298 297
rect 259 280 263 284
rect 289 282 293 286
rect 240 271 244 275
rect 339 293 343 297
rect 304 280 308 284
rect 334 282 338 286
rect 285 271 289 275
rect 384 293 388 297
rect 349 280 353 284
rect 379 282 383 286
rect 330 271 334 275
rect 429 293 433 297
rect 394 280 398 284
rect 424 282 428 286
rect 375 271 379 275
rect 474 293 478 297
rect 439 280 443 284
rect 469 282 473 286
rect 420 271 424 275
rect 519 293 523 297
rect 484 280 488 284
rect 514 282 518 286
rect 465 271 469 275
rect 564 293 568 297
rect 529 280 533 284
rect 559 282 563 286
rect 510 271 514 275
rect 609 293 613 297
rect 574 280 578 284
rect 604 282 608 286
rect 555 271 559 275
rect 654 293 658 297
rect 619 280 623 284
rect 649 282 653 286
rect 600 271 604 275
rect 699 293 703 297
rect 664 280 668 284
rect 694 282 698 286
rect 645 271 649 275
rect 744 293 748 297
rect 709 280 713 284
rect 739 282 743 286
rect 690 271 694 275
rect 789 293 793 297
rect 754 280 758 284
rect 784 282 788 286
rect 735 271 739 275
rect 834 293 838 297
rect 799 280 803 284
rect 829 282 833 286
rect 780 271 784 275
rect 879 293 883 297
rect 844 280 848 284
rect 874 282 878 286
rect 825 271 829 275
rect 889 280 893 284
rect 870 271 874 275
rect 24 248 28 252
rect 19 237 23 241
rect 69 248 73 252
rect 34 235 38 239
rect 64 237 68 241
rect 15 226 19 230
rect 114 248 118 252
rect 79 235 83 239
rect 109 237 113 241
rect 60 226 64 230
rect 159 248 163 252
rect 124 235 128 239
rect 154 237 158 241
rect 105 226 109 230
rect 204 248 208 252
rect 169 235 173 239
rect 199 237 203 241
rect 150 226 154 230
rect 249 248 253 252
rect 214 235 218 239
rect 244 237 248 241
rect 195 226 199 230
rect 294 248 298 252
rect 259 235 263 239
rect 289 237 293 241
rect 240 226 244 230
rect 339 248 343 252
rect 304 235 308 239
rect 334 237 338 241
rect 285 226 289 230
rect 384 248 388 252
rect 349 235 353 239
rect 379 237 383 241
rect 330 226 334 230
rect 429 248 433 252
rect 394 235 398 239
rect 424 237 428 241
rect 375 226 379 230
rect 474 248 478 252
rect 439 235 443 239
rect 469 237 473 241
rect 420 226 424 230
rect 519 248 523 252
rect 484 235 488 239
rect 514 237 518 241
rect 465 226 469 230
rect 564 248 568 252
rect 529 235 533 239
rect 559 237 563 241
rect 510 226 514 230
rect 609 248 613 252
rect 574 235 578 239
rect 604 237 608 241
rect 555 226 559 230
rect 654 248 658 252
rect 619 235 623 239
rect 649 237 653 241
rect 600 226 604 230
rect 699 248 703 252
rect 664 235 668 239
rect 694 237 698 241
rect 645 226 649 230
rect 744 248 748 252
rect 709 235 713 239
rect 739 237 743 241
rect 690 226 694 230
rect 789 248 793 252
rect 754 235 758 239
rect 784 237 788 241
rect 735 226 739 230
rect 834 248 838 252
rect 799 235 803 239
rect 829 237 833 241
rect 780 226 784 230
rect 879 248 883 252
rect 844 235 848 239
rect 874 237 878 241
rect 825 226 829 230
rect 889 235 893 239
rect 870 226 874 230
rect 24 203 28 207
rect 19 192 23 196
rect 69 203 73 207
rect 34 190 38 194
rect 64 192 68 196
rect 15 181 19 185
rect 114 203 118 207
rect 79 190 83 194
rect 109 192 113 196
rect 60 181 64 185
rect 159 203 163 207
rect 124 190 128 194
rect 154 192 158 196
rect 105 181 109 185
rect 204 203 208 207
rect 169 190 173 194
rect 199 192 203 196
rect 150 181 154 185
rect 249 203 253 207
rect 214 190 218 194
rect 244 192 248 196
rect 195 181 199 185
rect 294 203 298 207
rect 259 190 263 194
rect 289 192 293 196
rect 240 181 244 185
rect 339 203 343 207
rect 304 190 308 194
rect 334 192 338 196
rect 285 181 289 185
rect 384 203 388 207
rect 349 190 353 194
rect 379 192 383 196
rect 330 181 334 185
rect 429 203 433 207
rect 394 190 398 194
rect 424 192 428 196
rect 375 181 379 185
rect 474 203 478 207
rect 439 190 443 194
rect 469 192 473 196
rect 420 181 424 185
rect 519 203 523 207
rect 484 190 488 194
rect 514 192 518 196
rect 465 181 469 185
rect 564 203 568 207
rect 529 190 533 194
rect 559 192 563 196
rect 510 181 514 185
rect 609 203 613 207
rect 574 190 578 194
rect 604 192 608 196
rect 555 181 559 185
rect 654 203 658 207
rect 619 190 623 194
rect 649 192 653 196
rect 600 181 604 185
rect 699 203 703 207
rect 664 190 668 194
rect 694 192 698 196
rect 645 181 649 185
rect 744 203 748 207
rect 709 190 713 194
rect 739 192 743 196
rect 690 181 694 185
rect 789 203 793 207
rect 754 190 758 194
rect 784 192 788 196
rect 735 181 739 185
rect 834 203 838 207
rect 799 190 803 194
rect 829 192 833 196
rect 780 181 784 185
rect 879 203 883 207
rect 844 190 848 194
rect 874 192 878 196
rect 825 181 829 185
rect 889 190 893 194
rect 870 181 874 185
rect 24 158 28 162
rect 19 147 23 151
rect 69 158 73 162
rect 34 145 38 149
rect 64 147 68 151
rect 15 136 19 140
rect 114 158 118 162
rect 79 145 83 149
rect 109 147 113 151
rect 60 136 64 140
rect 159 158 163 162
rect 124 145 128 149
rect 154 147 158 151
rect 105 136 109 140
rect 204 158 208 162
rect 169 145 173 149
rect 199 147 203 151
rect 150 136 154 140
rect 249 158 253 162
rect 214 145 218 149
rect 244 147 248 151
rect 195 136 199 140
rect 294 158 298 162
rect 259 145 263 149
rect 289 147 293 151
rect 240 136 244 140
rect 339 158 343 162
rect 304 145 308 149
rect 334 147 338 151
rect 285 136 289 140
rect 384 158 388 162
rect 349 145 353 149
rect 379 147 383 151
rect 330 136 334 140
rect 429 158 433 162
rect 394 145 398 149
rect 424 147 428 151
rect 375 136 379 140
rect 474 158 478 162
rect 439 145 443 149
rect 469 147 473 151
rect 420 136 424 140
rect 519 158 523 162
rect 484 145 488 149
rect 514 147 518 151
rect 465 136 469 140
rect 564 158 568 162
rect 529 145 533 149
rect 559 147 563 151
rect 510 136 514 140
rect 609 158 613 162
rect 574 145 578 149
rect 604 147 608 151
rect 555 136 559 140
rect 654 158 658 162
rect 619 145 623 149
rect 649 147 653 151
rect 600 136 604 140
rect 699 158 703 162
rect 664 145 668 149
rect 694 147 698 151
rect 645 136 649 140
rect 744 158 748 162
rect 709 145 713 149
rect 739 147 743 151
rect 690 136 694 140
rect 789 158 793 162
rect 754 145 758 149
rect 784 147 788 151
rect 735 136 739 140
rect 834 158 838 162
rect 799 145 803 149
rect 829 147 833 151
rect 780 136 784 140
rect 879 158 883 162
rect 844 145 848 149
rect 874 147 878 151
rect 825 136 829 140
rect 889 145 893 149
rect 870 136 874 140
rect 24 113 28 117
rect 19 102 23 106
rect 69 113 73 117
rect 34 100 38 104
rect 64 102 68 106
rect 15 91 19 95
rect 114 113 118 117
rect 79 100 83 104
rect 109 102 113 106
rect 60 91 64 95
rect 159 113 163 117
rect 124 100 128 104
rect 154 102 158 106
rect 105 91 109 95
rect 204 113 208 117
rect 169 100 173 104
rect 199 102 203 106
rect 150 91 154 95
rect 249 113 253 117
rect 214 100 218 104
rect 244 102 248 106
rect 195 91 199 95
rect 294 113 298 117
rect 259 100 263 104
rect 289 102 293 106
rect 240 91 244 95
rect 339 113 343 117
rect 304 100 308 104
rect 334 102 338 106
rect 285 91 289 95
rect 384 113 388 117
rect 349 100 353 104
rect 379 102 383 106
rect 330 91 334 95
rect 429 113 433 117
rect 394 100 398 104
rect 424 102 428 106
rect 375 91 379 95
rect 474 113 478 117
rect 439 100 443 104
rect 469 102 473 106
rect 420 91 424 95
rect 519 113 523 117
rect 484 100 488 104
rect 514 102 518 106
rect 465 91 469 95
rect 564 113 568 117
rect 529 100 533 104
rect 559 102 563 106
rect 510 91 514 95
rect 609 113 613 117
rect 574 100 578 104
rect 604 102 608 106
rect 555 91 559 95
rect 654 113 658 117
rect 619 100 623 104
rect 649 102 653 106
rect 600 91 604 95
rect 699 113 703 117
rect 664 100 668 104
rect 694 102 698 106
rect 645 91 649 95
rect 744 113 748 117
rect 709 100 713 104
rect 739 102 743 106
rect 690 91 694 95
rect 789 113 793 117
rect 754 100 758 104
rect 784 102 788 106
rect 735 91 739 95
rect 834 113 838 117
rect 799 100 803 104
rect 829 102 833 106
rect 780 91 784 95
rect 879 113 883 117
rect 844 100 848 104
rect 874 102 878 106
rect 825 91 829 95
rect 889 100 893 104
rect 870 91 874 95
rect 24 68 28 72
rect 19 57 23 61
rect 69 68 73 72
rect 34 55 38 59
rect 64 57 68 61
rect 15 46 19 50
rect 114 68 118 72
rect 79 55 83 59
rect 109 57 113 61
rect 60 46 64 50
rect 159 68 163 72
rect 124 55 128 59
rect 154 57 158 61
rect 105 46 109 50
rect 204 68 208 72
rect 169 55 173 59
rect 199 57 203 61
rect 150 46 154 50
rect 249 68 253 72
rect 214 55 218 59
rect 244 57 248 61
rect 195 46 199 50
rect 294 68 298 72
rect 259 55 263 59
rect 289 57 293 61
rect 240 46 244 50
rect 339 68 343 72
rect 304 55 308 59
rect 334 57 338 61
rect 285 46 289 50
rect 384 68 388 72
rect 349 55 353 59
rect 379 57 383 61
rect 330 46 334 50
rect 429 68 433 72
rect 394 55 398 59
rect 424 57 428 61
rect 375 46 379 50
rect 474 68 478 72
rect 439 55 443 59
rect 469 57 473 61
rect 420 46 424 50
rect 519 68 523 72
rect 484 55 488 59
rect 514 57 518 61
rect 465 46 469 50
rect 564 68 568 72
rect 529 55 533 59
rect 559 57 563 61
rect 510 46 514 50
rect 609 68 613 72
rect 574 55 578 59
rect 604 57 608 61
rect 555 46 559 50
rect 654 68 658 72
rect 619 55 623 59
rect 649 57 653 61
rect 600 46 604 50
rect 699 68 703 72
rect 664 55 668 59
rect 694 57 698 61
rect 645 46 649 50
rect 744 68 748 72
rect 709 55 713 59
rect 739 57 743 61
rect 690 46 694 50
rect 789 68 793 72
rect 754 55 758 59
rect 784 57 788 61
rect 735 46 739 50
rect 834 68 838 72
rect 799 55 803 59
rect 829 57 833 61
rect 780 46 784 50
rect 879 68 883 72
rect 844 55 848 59
rect 874 57 878 61
rect 825 46 829 50
rect 889 55 893 59
rect 870 46 874 50
rect 24 23 28 27
rect 19 12 23 16
rect 69 23 73 27
rect 34 10 38 14
rect 64 12 68 16
rect 15 1 19 5
rect 114 23 118 27
rect 79 10 83 14
rect 109 12 113 16
rect 60 1 64 5
rect 159 23 163 27
rect 124 10 128 14
rect 154 12 158 16
rect 105 1 109 5
rect 204 23 208 27
rect 169 10 173 14
rect 199 12 203 16
rect 150 1 154 5
rect 249 23 253 27
rect 214 10 218 14
rect 244 12 248 16
rect 195 1 199 5
rect 294 23 298 27
rect 259 10 263 14
rect 289 12 293 16
rect 240 1 244 5
rect 339 23 343 27
rect 304 10 308 14
rect 334 12 338 16
rect 285 1 289 5
rect 384 23 388 27
rect 349 10 353 14
rect 379 12 383 16
rect 330 1 334 5
rect 429 23 433 27
rect 394 10 398 14
rect 424 12 428 16
rect 375 1 379 5
rect 474 23 478 27
rect 439 10 443 14
rect 469 12 473 16
rect 420 1 424 5
rect 519 23 523 27
rect 484 10 488 14
rect 514 12 518 16
rect 465 1 469 5
rect 564 23 568 27
rect 529 10 533 14
rect 559 12 563 16
rect 510 1 514 5
rect 609 23 613 27
rect 574 10 578 14
rect 604 12 608 16
rect 555 1 559 5
rect 654 23 658 27
rect 619 10 623 14
rect 649 12 653 16
rect 600 1 604 5
rect 699 23 703 27
rect 664 10 668 14
rect 694 12 698 16
rect 645 1 649 5
rect 744 23 748 27
rect 709 10 713 14
rect 739 12 743 16
rect 690 1 694 5
rect 789 23 793 27
rect 754 10 758 14
rect 784 12 788 16
rect 735 1 739 5
rect 834 23 838 27
rect 799 10 803 14
rect 829 12 833 16
rect 780 1 784 5
rect 879 23 883 27
rect 844 10 848 14
rect 874 12 878 16
rect 825 1 829 5
rect 889 10 893 14
rect 870 1 874 5
rect -296 -161 -292 -157
rect -273 -169 -269 -165
rect -192 -158 -188 -154
rect -197 -169 -193 -165
rect -286 -175 -282 -171
rect -182 -171 -178 -167
rect -201 -180 -197 -176
<< metal1 >>
rect 0 866 3 900
rect 35 875 38 900
rect 18 871 22 874
rect 31 872 38 875
rect 28 866 31 871
rect 0 863 8 866
rect 0 821 3 863
rect 28 858 31 862
rect 45 866 48 900
rect 80 875 83 900
rect 63 871 67 874
rect 76 872 83 875
rect 73 866 76 871
rect 45 863 53 866
rect 28 855 38 858
rect 35 830 38 855
rect 18 826 22 829
rect 31 827 38 830
rect 28 821 31 826
rect 0 818 8 821
rect 0 776 3 818
rect 28 813 31 817
rect 45 821 48 863
rect 73 858 76 862
rect 90 866 93 900
rect 125 875 128 900
rect 108 871 112 874
rect 121 872 128 875
rect 118 866 121 871
rect 90 863 98 866
rect 73 855 83 858
rect 80 830 83 855
rect 63 826 67 829
rect 76 827 83 830
rect 73 821 76 826
rect 45 818 53 821
rect 28 810 38 813
rect 35 785 38 810
rect 18 781 22 784
rect 31 782 38 785
rect 28 776 31 781
rect 0 773 8 776
rect 0 731 3 773
rect 28 768 31 772
rect 45 776 48 818
rect 73 813 76 817
rect 90 821 93 863
rect 118 858 121 862
rect 135 866 138 900
rect 170 875 173 900
rect 153 871 157 874
rect 166 872 173 875
rect 163 866 166 871
rect 135 863 143 866
rect 118 855 128 858
rect 125 830 128 855
rect 108 826 112 829
rect 121 827 128 830
rect 118 821 121 826
rect 90 818 98 821
rect 73 810 83 813
rect 80 785 83 810
rect 63 781 67 784
rect 76 782 83 785
rect 73 776 76 781
rect 45 773 53 776
rect 28 765 38 768
rect 35 740 38 765
rect 18 736 22 739
rect 31 737 38 740
rect 28 731 31 736
rect 0 728 8 731
rect 0 686 3 728
rect 28 723 31 727
rect 45 731 48 773
rect 73 768 76 772
rect 90 776 93 818
rect 118 813 121 817
rect 135 821 138 863
rect 163 858 166 862
rect 180 866 183 900
rect 215 875 218 900
rect 198 871 202 874
rect 211 872 218 875
rect 208 866 211 871
rect 180 863 188 866
rect 163 855 173 858
rect 170 830 173 855
rect 153 826 157 829
rect 166 827 173 830
rect 163 821 166 826
rect 135 818 143 821
rect 118 810 128 813
rect 125 785 128 810
rect 108 781 112 784
rect 121 782 128 785
rect 118 776 121 781
rect 90 773 98 776
rect 73 765 83 768
rect 80 740 83 765
rect 63 736 67 739
rect 76 737 83 740
rect 73 731 76 736
rect 45 728 53 731
rect 28 720 38 723
rect 35 695 38 720
rect 18 691 22 694
rect 31 692 38 695
rect 28 686 31 691
rect 0 683 8 686
rect 0 641 3 683
rect 28 678 31 682
rect 45 686 48 728
rect 73 723 76 727
rect 90 731 93 773
rect 118 768 121 772
rect 135 776 138 818
rect 163 813 166 817
rect 180 821 183 863
rect 208 858 211 862
rect 225 866 228 900
rect 260 875 263 900
rect 243 871 247 874
rect 256 872 263 875
rect 253 866 256 871
rect 225 863 233 866
rect 208 855 218 858
rect 215 830 218 855
rect 198 826 202 829
rect 211 827 218 830
rect 208 821 211 826
rect 180 818 188 821
rect 163 810 173 813
rect 170 785 173 810
rect 153 781 157 784
rect 166 782 173 785
rect 163 776 166 781
rect 135 773 143 776
rect 118 765 128 768
rect 125 740 128 765
rect 108 736 112 739
rect 121 737 128 740
rect 118 731 121 736
rect 90 728 98 731
rect 73 720 83 723
rect 80 695 83 720
rect 63 691 67 694
rect 76 692 83 695
rect 73 686 76 691
rect 45 683 53 686
rect 28 675 38 678
rect 35 650 38 675
rect 18 646 22 649
rect 31 647 38 650
rect 28 641 31 646
rect 0 638 8 641
rect 0 596 3 638
rect 28 633 31 637
rect 45 641 48 683
rect 73 678 76 682
rect 90 686 93 728
rect 118 723 121 727
rect 135 731 138 773
rect 163 768 166 772
rect 180 776 183 818
rect 208 813 211 817
rect 225 821 228 863
rect 253 858 256 862
rect 270 866 273 900
rect 305 875 308 900
rect 288 871 292 874
rect 301 872 308 875
rect 298 866 301 871
rect 270 863 278 866
rect 253 855 263 858
rect 260 830 263 855
rect 243 826 247 829
rect 256 827 263 830
rect 253 821 256 826
rect 225 818 233 821
rect 208 810 218 813
rect 215 785 218 810
rect 198 781 202 784
rect 211 782 218 785
rect 208 776 211 781
rect 180 773 188 776
rect 163 765 173 768
rect 170 740 173 765
rect 153 736 157 739
rect 166 737 173 740
rect 163 731 166 736
rect 135 728 143 731
rect 118 720 128 723
rect 125 695 128 720
rect 108 691 112 694
rect 121 692 128 695
rect 118 686 121 691
rect 90 683 98 686
rect 73 675 83 678
rect 80 650 83 675
rect 63 646 67 649
rect 76 647 83 650
rect 73 641 76 646
rect 45 638 53 641
rect 28 630 38 633
rect 35 605 38 630
rect 18 601 22 604
rect 31 602 38 605
rect 28 596 31 601
rect 0 593 8 596
rect 0 551 3 593
rect 28 588 31 592
rect 45 596 48 638
rect 73 633 76 637
rect 90 641 93 683
rect 118 678 121 682
rect 135 686 138 728
rect 163 723 166 727
rect 180 731 183 773
rect 208 768 211 772
rect 225 776 228 818
rect 253 813 256 817
rect 270 821 273 863
rect 298 858 301 862
rect 315 866 318 900
rect 350 875 353 900
rect 333 871 337 874
rect 346 872 353 875
rect 343 866 346 871
rect 315 863 323 866
rect 298 855 308 858
rect 305 830 308 855
rect 288 826 292 829
rect 301 827 308 830
rect 298 821 301 826
rect 270 818 278 821
rect 253 810 263 813
rect 260 785 263 810
rect 243 781 247 784
rect 256 782 263 785
rect 253 776 256 781
rect 225 773 233 776
rect 208 765 218 768
rect 215 740 218 765
rect 198 736 202 739
rect 211 737 218 740
rect 208 731 211 736
rect 180 728 188 731
rect 163 720 173 723
rect 170 695 173 720
rect 153 691 157 694
rect 166 692 173 695
rect 163 686 166 691
rect 135 683 143 686
rect 118 675 128 678
rect 125 650 128 675
rect 108 646 112 649
rect 121 647 128 650
rect 118 641 121 646
rect 90 638 98 641
rect 73 630 83 633
rect 80 605 83 630
rect 63 601 67 604
rect 76 602 83 605
rect 73 596 76 601
rect 45 593 53 596
rect 28 585 38 588
rect 35 560 38 585
rect 18 556 22 559
rect 31 557 38 560
rect 28 551 31 556
rect 0 548 8 551
rect 0 506 3 548
rect 28 543 31 547
rect 45 551 48 593
rect 73 588 76 592
rect 90 596 93 638
rect 118 633 121 637
rect 135 641 138 683
rect 163 678 166 682
rect 180 686 183 728
rect 208 723 211 727
rect 225 731 228 773
rect 253 768 256 772
rect 270 776 273 818
rect 298 813 301 817
rect 315 821 318 863
rect 343 858 346 862
rect 360 866 363 900
rect 395 875 398 900
rect 378 871 382 874
rect 391 872 398 875
rect 388 866 391 871
rect 360 863 368 866
rect 343 855 353 858
rect 350 830 353 855
rect 333 826 337 829
rect 346 827 353 830
rect 343 821 346 826
rect 315 818 323 821
rect 298 810 308 813
rect 305 785 308 810
rect 288 781 292 784
rect 301 782 308 785
rect 298 776 301 781
rect 270 773 278 776
rect 253 765 263 768
rect 260 740 263 765
rect 243 736 247 739
rect 256 737 263 740
rect 253 731 256 736
rect 225 728 233 731
rect 208 720 218 723
rect 215 695 218 720
rect 198 691 202 694
rect 211 692 218 695
rect 208 686 211 691
rect 180 683 188 686
rect 163 675 173 678
rect 170 650 173 675
rect 153 646 157 649
rect 166 647 173 650
rect 163 641 166 646
rect 135 638 143 641
rect 118 630 128 633
rect 125 605 128 630
rect 108 601 112 604
rect 121 602 128 605
rect 118 596 121 601
rect 90 593 98 596
rect 73 585 83 588
rect 80 560 83 585
rect 63 556 67 559
rect 76 557 83 560
rect 73 551 76 556
rect 45 548 53 551
rect 28 540 38 543
rect 35 515 38 540
rect 18 511 22 514
rect 31 512 38 515
rect 28 506 31 511
rect 0 503 8 506
rect 0 461 3 503
rect 28 498 31 502
rect 45 506 48 548
rect 73 543 76 547
rect 90 551 93 593
rect 118 588 121 592
rect 135 596 138 638
rect 163 633 166 637
rect 180 641 183 683
rect 208 678 211 682
rect 225 686 228 728
rect 253 723 256 727
rect 270 731 273 773
rect 298 768 301 772
rect 315 776 318 818
rect 343 813 346 817
rect 360 821 363 863
rect 388 858 391 862
rect 405 866 408 900
rect 440 875 443 900
rect 423 871 427 874
rect 436 872 443 875
rect 433 866 436 871
rect 405 863 413 866
rect 388 855 398 858
rect 395 830 398 855
rect 378 826 382 829
rect 391 827 398 830
rect 388 821 391 826
rect 360 818 368 821
rect 343 810 353 813
rect 350 785 353 810
rect 333 781 337 784
rect 346 782 353 785
rect 343 776 346 781
rect 315 773 323 776
rect 298 765 308 768
rect 305 740 308 765
rect 288 736 292 739
rect 301 737 308 740
rect 298 731 301 736
rect 270 728 278 731
rect 253 720 263 723
rect 260 695 263 720
rect 243 691 247 694
rect 256 692 263 695
rect 253 686 256 691
rect 225 683 233 686
rect 208 675 218 678
rect 215 650 218 675
rect 198 646 202 649
rect 211 647 218 650
rect 208 641 211 646
rect 180 638 188 641
rect 163 630 173 633
rect 170 605 173 630
rect 153 601 157 604
rect 166 602 173 605
rect 163 596 166 601
rect 135 593 143 596
rect 118 585 128 588
rect 125 560 128 585
rect 108 556 112 559
rect 121 557 128 560
rect 118 551 121 556
rect 90 548 98 551
rect 73 540 83 543
rect 80 515 83 540
rect 63 511 67 514
rect 76 512 83 515
rect 73 506 76 511
rect 45 503 53 506
rect 28 495 38 498
rect 35 470 38 495
rect 18 466 22 469
rect 31 467 38 470
rect 28 461 31 466
rect 0 458 8 461
rect 0 416 3 458
rect 28 453 31 457
rect 45 461 48 503
rect 73 498 76 502
rect 90 506 93 548
rect 118 543 121 547
rect 135 551 138 593
rect 163 588 166 592
rect 180 596 183 638
rect 208 633 211 637
rect 225 641 228 683
rect 253 678 256 682
rect 270 686 273 728
rect 298 723 301 727
rect 315 731 318 773
rect 343 768 346 772
rect 360 776 363 818
rect 388 813 391 817
rect 405 821 408 863
rect 433 858 436 862
rect 450 866 453 900
rect 485 875 488 900
rect 468 871 472 874
rect 481 872 488 875
rect 478 866 481 871
rect 450 863 458 866
rect 433 855 443 858
rect 440 830 443 855
rect 423 826 427 829
rect 436 827 443 830
rect 433 821 436 826
rect 405 818 413 821
rect 388 810 398 813
rect 395 785 398 810
rect 378 781 382 784
rect 391 782 398 785
rect 388 776 391 781
rect 360 773 368 776
rect 343 765 353 768
rect 350 740 353 765
rect 333 736 337 739
rect 346 737 353 740
rect 343 731 346 736
rect 315 728 323 731
rect 298 720 308 723
rect 305 695 308 720
rect 288 691 292 694
rect 301 692 308 695
rect 298 686 301 691
rect 270 683 278 686
rect 253 675 263 678
rect 260 650 263 675
rect 243 646 247 649
rect 256 647 263 650
rect 253 641 256 646
rect 225 638 233 641
rect 208 630 218 633
rect 215 605 218 630
rect 198 601 202 604
rect 211 602 218 605
rect 208 596 211 601
rect 180 593 188 596
rect 163 585 173 588
rect 170 560 173 585
rect 153 556 157 559
rect 166 557 173 560
rect 163 551 166 556
rect 135 548 143 551
rect 118 540 128 543
rect 125 515 128 540
rect 108 511 112 514
rect 121 512 128 515
rect 118 506 121 511
rect 90 503 98 506
rect 73 495 83 498
rect 80 470 83 495
rect 63 466 67 469
rect 76 467 83 470
rect 73 461 76 466
rect 45 458 53 461
rect 28 450 38 453
rect 35 425 38 450
rect 18 421 22 424
rect 31 422 38 425
rect 28 416 31 421
rect 0 413 8 416
rect 0 371 3 413
rect 28 408 31 412
rect 45 416 48 458
rect 73 453 76 457
rect 90 461 93 503
rect 118 498 121 502
rect 135 506 138 548
rect 163 543 166 547
rect 180 551 183 593
rect 208 588 211 592
rect 225 596 228 638
rect 253 633 256 637
rect 270 641 273 683
rect 298 678 301 682
rect 315 686 318 728
rect 343 723 346 727
rect 360 731 363 773
rect 388 768 391 772
rect 405 776 408 818
rect 433 813 436 817
rect 450 821 453 863
rect 478 858 481 862
rect 495 866 498 900
rect 530 875 533 900
rect 513 871 517 874
rect 526 872 533 875
rect 523 866 526 871
rect 495 863 503 866
rect 478 855 488 858
rect 485 830 488 855
rect 468 826 472 829
rect 481 827 488 830
rect 478 821 481 826
rect 450 818 458 821
rect 433 810 443 813
rect 440 785 443 810
rect 423 781 427 784
rect 436 782 443 785
rect 433 776 436 781
rect 405 773 413 776
rect 388 765 398 768
rect 395 740 398 765
rect 378 736 382 739
rect 391 737 398 740
rect 388 731 391 736
rect 360 728 368 731
rect 343 720 353 723
rect 350 695 353 720
rect 333 691 337 694
rect 346 692 353 695
rect 343 686 346 691
rect 315 683 323 686
rect 298 675 308 678
rect 305 650 308 675
rect 288 646 292 649
rect 301 647 308 650
rect 298 641 301 646
rect 270 638 278 641
rect 253 630 263 633
rect 260 605 263 630
rect 243 601 247 604
rect 256 602 263 605
rect 253 596 256 601
rect 225 593 233 596
rect 208 585 218 588
rect 215 560 218 585
rect 198 556 202 559
rect 211 557 218 560
rect 208 551 211 556
rect 180 548 188 551
rect 163 540 173 543
rect 170 515 173 540
rect 153 511 157 514
rect 166 512 173 515
rect 163 506 166 511
rect 135 503 143 506
rect 118 495 128 498
rect 125 470 128 495
rect 108 466 112 469
rect 121 467 128 470
rect 118 461 121 466
rect 90 458 98 461
rect 73 450 83 453
rect 80 425 83 450
rect 63 421 67 424
rect 76 422 83 425
rect 73 416 76 421
rect 45 413 53 416
rect 28 405 38 408
rect 35 380 38 405
rect 18 376 22 379
rect 31 377 38 380
rect 28 371 31 376
rect 0 368 8 371
rect 0 326 3 368
rect 28 363 31 367
rect 45 371 48 413
rect 73 408 76 412
rect 90 416 93 458
rect 118 453 121 457
rect 135 461 138 503
rect 163 498 166 502
rect 180 506 183 548
rect 208 543 211 547
rect 225 551 228 593
rect 253 588 256 592
rect 270 596 273 638
rect 298 633 301 637
rect 315 641 318 683
rect 343 678 346 682
rect 360 686 363 728
rect 388 723 391 727
rect 405 731 408 773
rect 433 768 436 772
rect 450 776 453 818
rect 478 813 481 817
rect 495 821 498 863
rect 523 858 526 862
rect 540 866 543 900
rect 575 875 578 900
rect 558 871 562 874
rect 571 872 578 875
rect 568 866 571 871
rect 540 863 548 866
rect 523 855 533 858
rect 530 830 533 855
rect 513 826 517 829
rect 526 827 533 830
rect 523 821 526 826
rect 495 818 503 821
rect 478 810 488 813
rect 485 785 488 810
rect 468 781 472 784
rect 481 782 488 785
rect 478 776 481 781
rect 450 773 458 776
rect 433 765 443 768
rect 440 740 443 765
rect 423 736 427 739
rect 436 737 443 740
rect 433 731 436 736
rect 405 728 413 731
rect 388 720 398 723
rect 395 695 398 720
rect 378 691 382 694
rect 391 692 398 695
rect 388 686 391 691
rect 360 683 368 686
rect 343 675 353 678
rect 350 650 353 675
rect 333 646 337 649
rect 346 647 353 650
rect 343 641 346 646
rect 315 638 323 641
rect 298 630 308 633
rect 305 605 308 630
rect 288 601 292 604
rect 301 602 308 605
rect 298 596 301 601
rect 270 593 278 596
rect 253 585 263 588
rect 260 560 263 585
rect 243 556 247 559
rect 256 557 263 560
rect 253 551 256 556
rect 225 548 233 551
rect 208 540 218 543
rect 215 515 218 540
rect 198 511 202 514
rect 211 512 218 515
rect 208 506 211 511
rect 180 503 188 506
rect 163 495 173 498
rect 170 470 173 495
rect 153 466 157 469
rect 166 467 173 470
rect 163 461 166 466
rect 135 458 143 461
rect 118 450 128 453
rect 125 425 128 450
rect 108 421 112 424
rect 121 422 128 425
rect 118 416 121 421
rect 90 413 98 416
rect 73 405 83 408
rect 80 380 83 405
rect 63 376 67 379
rect 76 377 83 380
rect 73 371 76 376
rect 45 368 53 371
rect 28 360 38 363
rect 35 335 38 360
rect 18 331 22 334
rect 31 332 38 335
rect 28 326 31 331
rect 0 323 8 326
rect 0 281 3 323
rect 28 318 31 322
rect 45 326 48 368
rect 73 363 76 367
rect 90 371 93 413
rect 118 408 121 412
rect 135 416 138 458
rect 163 453 166 457
rect 180 461 183 503
rect 208 498 211 502
rect 225 506 228 548
rect 253 543 256 547
rect 270 551 273 593
rect 298 588 301 592
rect 315 596 318 638
rect 343 633 346 637
rect 360 641 363 683
rect 388 678 391 682
rect 405 686 408 728
rect 433 723 436 727
rect 450 731 453 773
rect 478 768 481 772
rect 495 776 498 818
rect 523 813 526 817
rect 540 821 543 863
rect 568 858 571 862
rect 585 866 588 900
rect 620 875 623 900
rect 603 871 607 874
rect 616 872 623 875
rect 613 866 616 871
rect 585 863 593 866
rect 568 855 578 858
rect 575 830 578 855
rect 558 826 562 829
rect 571 827 578 830
rect 568 821 571 826
rect 540 818 548 821
rect 523 810 533 813
rect 530 785 533 810
rect 513 781 517 784
rect 526 782 533 785
rect 523 776 526 781
rect 495 773 503 776
rect 478 765 488 768
rect 485 740 488 765
rect 468 736 472 739
rect 481 737 488 740
rect 478 731 481 736
rect 450 728 458 731
rect 433 720 443 723
rect 440 695 443 720
rect 423 691 427 694
rect 436 692 443 695
rect 433 686 436 691
rect 405 683 413 686
rect 388 675 398 678
rect 395 650 398 675
rect 378 646 382 649
rect 391 647 398 650
rect 388 641 391 646
rect 360 638 368 641
rect 343 630 353 633
rect 350 605 353 630
rect 333 601 337 604
rect 346 602 353 605
rect 343 596 346 601
rect 315 593 323 596
rect 298 585 308 588
rect 305 560 308 585
rect 288 556 292 559
rect 301 557 308 560
rect 298 551 301 556
rect 270 548 278 551
rect 253 540 263 543
rect 260 515 263 540
rect 243 511 247 514
rect 256 512 263 515
rect 253 506 256 511
rect 225 503 233 506
rect 208 495 218 498
rect 215 470 218 495
rect 198 466 202 469
rect 211 467 218 470
rect 208 461 211 466
rect 180 458 188 461
rect 163 450 173 453
rect 170 425 173 450
rect 153 421 157 424
rect 166 422 173 425
rect 163 416 166 421
rect 135 413 143 416
rect 118 405 128 408
rect 125 380 128 405
rect 108 376 112 379
rect 121 377 128 380
rect 118 371 121 376
rect 90 368 98 371
rect 73 360 83 363
rect 80 335 83 360
rect 63 331 67 334
rect 76 332 83 335
rect 73 326 76 331
rect 45 323 53 326
rect 28 315 38 318
rect 35 290 38 315
rect 18 286 22 289
rect 31 287 38 290
rect 28 281 31 286
rect 0 278 8 281
rect 0 236 3 278
rect 28 273 31 277
rect 45 281 48 323
rect 73 318 76 322
rect 90 326 93 368
rect 118 363 121 367
rect 135 371 138 413
rect 163 408 166 412
rect 180 416 183 458
rect 208 453 211 457
rect 225 461 228 503
rect 253 498 256 502
rect 270 506 273 548
rect 298 543 301 547
rect 315 551 318 593
rect 343 588 346 592
rect 360 596 363 638
rect 388 633 391 637
rect 405 641 408 683
rect 433 678 436 682
rect 450 686 453 728
rect 478 723 481 727
rect 495 731 498 773
rect 523 768 526 772
rect 540 776 543 818
rect 568 813 571 817
rect 585 821 588 863
rect 613 858 616 862
rect 630 866 633 900
rect 665 875 668 900
rect 648 871 652 874
rect 661 872 668 875
rect 658 866 661 871
rect 630 863 638 866
rect 613 855 623 858
rect 620 830 623 855
rect 603 826 607 829
rect 616 827 623 830
rect 613 821 616 826
rect 585 818 593 821
rect 568 810 578 813
rect 575 785 578 810
rect 558 781 562 784
rect 571 782 578 785
rect 568 776 571 781
rect 540 773 548 776
rect 523 765 533 768
rect 530 740 533 765
rect 513 736 517 739
rect 526 737 533 740
rect 523 731 526 736
rect 495 728 503 731
rect 478 720 488 723
rect 485 695 488 720
rect 468 691 472 694
rect 481 692 488 695
rect 478 686 481 691
rect 450 683 458 686
rect 433 675 443 678
rect 440 650 443 675
rect 423 646 427 649
rect 436 647 443 650
rect 433 641 436 646
rect 405 638 413 641
rect 388 630 398 633
rect 395 605 398 630
rect 378 601 382 604
rect 391 602 398 605
rect 388 596 391 601
rect 360 593 368 596
rect 343 585 353 588
rect 350 560 353 585
rect 333 556 337 559
rect 346 557 353 560
rect 343 551 346 556
rect 315 548 323 551
rect 298 540 308 543
rect 305 515 308 540
rect 288 511 292 514
rect 301 512 308 515
rect 298 506 301 511
rect 270 503 278 506
rect 253 495 263 498
rect 260 470 263 495
rect 243 466 247 469
rect 256 467 263 470
rect 253 461 256 466
rect 225 458 233 461
rect 208 450 218 453
rect 215 425 218 450
rect 198 421 202 424
rect 211 422 218 425
rect 208 416 211 421
rect 180 413 188 416
rect 163 405 173 408
rect 170 380 173 405
rect 153 376 157 379
rect 166 377 173 380
rect 163 371 166 376
rect 135 368 143 371
rect 118 360 128 363
rect 125 335 128 360
rect 108 331 112 334
rect 121 332 128 335
rect 118 326 121 331
rect 90 323 98 326
rect 73 315 83 318
rect 80 290 83 315
rect 63 286 67 289
rect 76 287 83 290
rect 73 281 76 286
rect 45 278 53 281
rect 28 270 38 273
rect 35 245 38 270
rect 18 241 22 244
rect 31 242 38 245
rect 28 236 31 241
rect 0 233 8 236
rect 0 191 3 233
rect 28 228 31 232
rect 45 236 48 278
rect 73 273 76 277
rect 90 281 93 323
rect 118 318 121 322
rect 135 326 138 368
rect 163 363 166 367
rect 180 371 183 413
rect 208 408 211 412
rect 225 416 228 458
rect 253 453 256 457
rect 270 461 273 503
rect 298 498 301 502
rect 315 506 318 548
rect 343 543 346 547
rect 360 551 363 593
rect 388 588 391 592
rect 405 596 408 638
rect 433 633 436 637
rect 450 641 453 683
rect 478 678 481 682
rect 495 686 498 728
rect 523 723 526 727
rect 540 731 543 773
rect 568 768 571 772
rect 585 776 588 818
rect 613 813 616 817
rect 630 821 633 863
rect 658 858 661 862
rect 675 866 678 900
rect 710 875 713 900
rect 693 871 697 874
rect 706 872 713 875
rect 703 866 706 871
rect 675 863 683 866
rect 658 855 668 858
rect 665 830 668 855
rect 648 826 652 829
rect 661 827 668 830
rect 658 821 661 826
rect 630 818 638 821
rect 613 810 623 813
rect 620 785 623 810
rect 603 781 607 784
rect 616 782 623 785
rect 613 776 616 781
rect 585 773 593 776
rect 568 765 578 768
rect 575 740 578 765
rect 558 736 562 739
rect 571 737 578 740
rect 568 731 571 736
rect 540 728 548 731
rect 523 720 533 723
rect 530 695 533 720
rect 513 691 517 694
rect 526 692 533 695
rect 523 686 526 691
rect 495 683 503 686
rect 478 675 488 678
rect 485 650 488 675
rect 468 646 472 649
rect 481 647 488 650
rect 478 641 481 646
rect 450 638 458 641
rect 433 630 443 633
rect 440 605 443 630
rect 423 601 427 604
rect 436 602 443 605
rect 433 596 436 601
rect 405 593 413 596
rect 388 585 398 588
rect 395 560 398 585
rect 378 556 382 559
rect 391 557 398 560
rect 388 551 391 556
rect 360 548 368 551
rect 343 540 353 543
rect 350 515 353 540
rect 333 511 337 514
rect 346 512 353 515
rect 343 506 346 511
rect 315 503 323 506
rect 298 495 308 498
rect 305 470 308 495
rect 288 466 292 469
rect 301 467 308 470
rect 298 461 301 466
rect 270 458 278 461
rect 253 450 263 453
rect 260 425 263 450
rect 243 421 247 424
rect 256 422 263 425
rect 253 416 256 421
rect 225 413 233 416
rect 208 405 218 408
rect 215 380 218 405
rect 198 376 202 379
rect 211 377 218 380
rect 208 371 211 376
rect 180 368 188 371
rect 163 360 173 363
rect 170 335 173 360
rect 153 331 157 334
rect 166 332 173 335
rect 163 326 166 331
rect 135 323 143 326
rect 118 315 128 318
rect 125 290 128 315
rect 108 286 112 289
rect 121 287 128 290
rect 118 281 121 286
rect 90 278 98 281
rect 73 270 83 273
rect 80 245 83 270
rect 63 241 67 244
rect 76 242 83 245
rect 73 236 76 241
rect 45 233 53 236
rect 28 225 38 228
rect 35 200 38 225
rect 18 196 22 199
rect 31 197 38 200
rect 28 191 31 196
rect 0 188 8 191
rect 0 146 3 188
rect 28 183 31 187
rect 45 191 48 233
rect 73 228 76 232
rect 90 236 93 278
rect 118 273 121 277
rect 135 281 138 323
rect 163 318 166 322
rect 180 326 183 368
rect 208 363 211 367
rect 225 371 228 413
rect 253 408 256 412
rect 270 416 273 458
rect 298 453 301 457
rect 315 461 318 503
rect 343 498 346 502
rect 360 506 363 548
rect 388 543 391 547
rect 405 551 408 593
rect 433 588 436 592
rect 450 596 453 638
rect 478 633 481 637
rect 495 641 498 683
rect 523 678 526 682
rect 540 686 543 728
rect 568 723 571 727
rect 585 731 588 773
rect 613 768 616 772
rect 630 776 633 818
rect 658 813 661 817
rect 675 821 678 863
rect 703 858 706 862
rect 720 866 723 900
rect 755 875 758 900
rect 738 871 742 874
rect 751 872 758 875
rect 748 866 751 871
rect 720 863 728 866
rect 703 855 713 858
rect 710 830 713 855
rect 693 826 697 829
rect 706 827 713 830
rect 703 821 706 826
rect 675 818 683 821
rect 658 810 668 813
rect 665 785 668 810
rect 648 781 652 784
rect 661 782 668 785
rect 658 776 661 781
rect 630 773 638 776
rect 613 765 623 768
rect 620 740 623 765
rect 603 736 607 739
rect 616 737 623 740
rect 613 731 616 736
rect 585 728 593 731
rect 568 720 578 723
rect 575 695 578 720
rect 558 691 562 694
rect 571 692 578 695
rect 568 686 571 691
rect 540 683 548 686
rect 523 675 533 678
rect 530 650 533 675
rect 513 646 517 649
rect 526 647 533 650
rect 523 641 526 646
rect 495 638 503 641
rect 478 630 488 633
rect 485 605 488 630
rect 468 601 472 604
rect 481 602 488 605
rect 478 596 481 601
rect 450 593 458 596
rect 433 585 443 588
rect 440 560 443 585
rect 423 556 427 559
rect 436 557 443 560
rect 433 551 436 556
rect 405 548 413 551
rect 388 540 398 543
rect 395 515 398 540
rect 378 511 382 514
rect 391 512 398 515
rect 388 506 391 511
rect 360 503 368 506
rect 343 495 353 498
rect 350 470 353 495
rect 333 466 337 469
rect 346 467 353 470
rect 343 461 346 466
rect 315 458 323 461
rect 298 450 308 453
rect 305 425 308 450
rect 288 421 292 424
rect 301 422 308 425
rect 298 416 301 421
rect 270 413 278 416
rect 253 405 263 408
rect 260 380 263 405
rect 243 376 247 379
rect 256 377 263 380
rect 253 371 256 376
rect 225 368 233 371
rect 208 360 218 363
rect 215 335 218 360
rect 198 331 202 334
rect 211 332 218 335
rect 208 326 211 331
rect 180 323 188 326
rect 163 315 173 318
rect 170 290 173 315
rect 153 286 157 289
rect 166 287 173 290
rect 163 281 166 286
rect 135 278 143 281
rect 118 270 128 273
rect 125 245 128 270
rect 108 241 112 244
rect 121 242 128 245
rect 118 236 121 241
rect 90 233 98 236
rect 73 225 83 228
rect 80 200 83 225
rect 63 196 67 199
rect 76 197 83 200
rect 73 191 76 196
rect 45 188 53 191
rect 28 180 38 183
rect 35 155 38 180
rect 18 151 22 154
rect 31 152 38 155
rect 28 146 31 151
rect 0 143 8 146
rect 0 101 3 143
rect 28 138 31 142
rect 45 146 48 188
rect 73 183 76 187
rect 90 191 93 233
rect 118 228 121 232
rect 135 236 138 278
rect 163 273 166 277
rect 180 281 183 323
rect 208 318 211 322
rect 225 326 228 368
rect 253 363 256 367
rect 270 371 273 413
rect 298 408 301 412
rect 315 416 318 458
rect 343 453 346 457
rect 360 461 363 503
rect 388 498 391 502
rect 405 506 408 548
rect 433 543 436 547
rect 450 551 453 593
rect 478 588 481 592
rect 495 596 498 638
rect 523 633 526 637
rect 540 641 543 683
rect 568 678 571 682
rect 585 686 588 728
rect 613 723 616 727
rect 630 731 633 773
rect 658 768 661 772
rect 675 776 678 818
rect 703 813 706 817
rect 720 821 723 863
rect 748 858 751 862
rect 765 866 768 900
rect 800 875 803 900
rect 783 871 787 874
rect 796 872 803 875
rect 793 866 796 871
rect 765 863 773 866
rect 748 855 758 858
rect 755 830 758 855
rect 738 826 742 829
rect 751 827 758 830
rect 748 821 751 826
rect 720 818 728 821
rect 703 810 713 813
rect 710 785 713 810
rect 693 781 697 784
rect 706 782 713 785
rect 703 776 706 781
rect 675 773 683 776
rect 658 765 668 768
rect 665 740 668 765
rect 648 736 652 739
rect 661 737 668 740
rect 658 731 661 736
rect 630 728 638 731
rect 613 720 623 723
rect 620 695 623 720
rect 603 691 607 694
rect 616 692 623 695
rect 613 686 616 691
rect 585 683 593 686
rect 568 675 578 678
rect 575 650 578 675
rect 558 646 562 649
rect 571 647 578 650
rect 568 641 571 646
rect 540 638 548 641
rect 523 630 533 633
rect 530 605 533 630
rect 513 601 517 604
rect 526 602 533 605
rect 523 596 526 601
rect 495 593 503 596
rect 478 585 488 588
rect 485 560 488 585
rect 468 556 472 559
rect 481 557 488 560
rect 478 551 481 556
rect 450 548 458 551
rect 433 540 443 543
rect 440 515 443 540
rect 423 511 427 514
rect 436 512 443 515
rect 433 506 436 511
rect 405 503 413 506
rect 388 495 398 498
rect 395 470 398 495
rect 378 466 382 469
rect 391 467 398 470
rect 388 461 391 466
rect 360 458 368 461
rect 343 450 353 453
rect 350 425 353 450
rect 333 421 337 424
rect 346 422 353 425
rect 343 416 346 421
rect 315 413 323 416
rect 298 405 308 408
rect 305 380 308 405
rect 288 376 292 379
rect 301 377 308 380
rect 298 371 301 376
rect 270 368 278 371
rect 253 360 263 363
rect 260 335 263 360
rect 243 331 247 334
rect 256 332 263 335
rect 253 326 256 331
rect 225 323 233 326
rect 208 315 218 318
rect 215 290 218 315
rect 198 286 202 289
rect 211 287 218 290
rect 208 281 211 286
rect 180 278 188 281
rect 163 270 173 273
rect 170 245 173 270
rect 153 241 157 244
rect 166 242 173 245
rect 163 236 166 241
rect 135 233 143 236
rect 118 225 128 228
rect 125 200 128 225
rect 108 196 112 199
rect 121 197 128 200
rect 118 191 121 196
rect 90 188 98 191
rect 73 180 83 183
rect 80 155 83 180
rect 63 151 67 154
rect 76 152 83 155
rect 73 146 76 151
rect 45 143 53 146
rect 28 135 38 138
rect 35 110 38 135
rect 18 106 22 109
rect 31 107 38 110
rect 28 101 31 106
rect 0 98 8 101
rect 0 56 3 98
rect 28 93 31 97
rect 45 101 48 143
rect 73 138 76 142
rect 90 146 93 188
rect 118 183 121 187
rect 135 191 138 233
rect 163 228 166 232
rect 180 236 183 278
rect 208 273 211 277
rect 225 281 228 323
rect 253 318 256 322
rect 270 326 273 368
rect 298 363 301 367
rect 315 371 318 413
rect 343 408 346 412
rect 360 416 363 458
rect 388 453 391 457
rect 405 461 408 503
rect 433 498 436 502
rect 450 506 453 548
rect 478 543 481 547
rect 495 551 498 593
rect 523 588 526 592
rect 540 596 543 638
rect 568 633 571 637
rect 585 641 588 683
rect 613 678 616 682
rect 630 686 633 728
rect 658 723 661 727
rect 675 731 678 773
rect 703 768 706 772
rect 720 776 723 818
rect 748 813 751 817
rect 765 821 768 863
rect 793 858 796 862
rect 810 866 813 900
rect 845 875 848 900
rect 828 871 832 874
rect 841 872 848 875
rect 838 866 841 871
rect 810 863 818 866
rect 793 855 803 858
rect 800 830 803 855
rect 783 826 787 829
rect 796 827 803 830
rect 793 821 796 826
rect 765 818 773 821
rect 748 810 758 813
rect 755 785 758 810
rect 738 781 742 784
rect 751 782 758 785
rect 748 776 751 781
rect 720 773 728 776
rect 703 765 713 768
rect 710 740 713 765
rect 693 736 697 739
rect 706 737 713 740
rect 703 731 706 736
rect 675 728 683 731
rect 658 720 668 723
rect 665 695 668 720
rect 648 691 652 694
rect 661 692 668 695
rect 658 686 661 691
rect 630 683 638 686
rect 613 675 623 678
rect 620 650 623 675
rect 603 646 607 649
rect 616 647 623 650
rect 613 641 616 646
rect 585 638 593 641
rect 568 630 578 633
rect 575 605 578 630
rect 558 601 562 604
rect 571 602 578 605
rect 568 596 571 601
rect 540 593 548 596
rect 523 585 533 588
rect 530 560 533 585
rect 513 556 517 559
rect 526 557 533 560
rect 523 551 526 556
rect 495 548 503 551
rect 478 540 488 543
rect 485 515 488 540
rect 468 511 472 514
rect 481 512 488 515
rect 478 506 481 511
rect 450 503 458 506
rect 433 495 443 498
rect 440 470 443 495
rect 423 466 427 469
rect 436 467 443 470
rect 433 461 436 466
rect 405 458 413 461
rect 388 450 398 453
rect 395 425 398 450
rect 378 421 382 424
rect 391 422 398 425
rect 388 416 391 421
rect 360 413 368 416
rect 343 405 353 408
rect 350 380 353 405
rect 333 376 337 379
rect 346 377 353 380
rect 343 371 346 376
rect 315 368 323 371
rect 298 360 308 363
rect 305 335 308 360
rect 288 331 292 334
rect 301 332 308 335
rect 298 326 301 331
rect 270 323 278 326
rect 253 315 263 318
rect 260 290 263 315
rect 243 286 247 289
rect 256 287 263 290
rect 253 281 256 286
rect 225 278 233 281
rect 208 270 218 273
rect 215 245 218 270
rect 198 241 202 244
rect 211 242 218 245
rect 208 236 211 241
rect 180 233 188 236
rect 163 225 173 228
rect 170 200 173 225
rect 153 196 157 199
rect 166 197 173 200
rect 163 191 166 196
rect 135 188 143 191
rect 118 180 128 183
rect 125 155 128 180
rect 108 151 112 154
rect 121 152 128 155
rect 118 146 121 151
rect 90 143 98 146
rect 73 135 83 138
rect 80 110 83 135
rect 63 106 67 109
rect 76 107 83 110
rect 73 101 76 106
rect 45 98 53 101
rect 28 90 38 93
rect 35 65 38 90
rect 18 61 22 64
rect 31 62 38 65
rect 28 56 31 61
rect 0 53 8 56
rect 0 11 3 53
rect 28 48 31 52
rect 45 56 48 98
rect 73 93 76 97
rect 90 101 93 143
rect 118 138 121 142
rect 135 146 138 188
rect 163 183 166 187
rect 180 191 183 233
rect 208 228 211 232
rect 225 236 228 278
rect 253 273 256 277
rect 270 281 273 323
rect 298 318 301 322
rect 315 326 318 368
rect 343 363 346 367
rect 360 371 363 413
rect 388 408 391 412
rect 405 416 408 458
rect 433 453 436 457
rect 450 461 453 503
rect 478 498 481 502
rect 495 506 498 548
rect 523 543 526 547
rect 540 551 543 593
rect 568 588 571 592
rect 585 596 588 638
rect 613 633 616 637
rect 630 641 633 683
rect 658 678 661 682
rect 675 686 678 728
rect 703 723 706 727
rect 720 731 723 773
rect 748 768 751 772
rect 765 776 768 818
rect 793 813 796 817
rect 810 821 813 863
rect 838 858 841 862
rect 855 866 858 900
rect 890 875 893 900
rect 873 871 877 874
rect 886 872 893 875
rect 883 866 886 871
rect 855 863 863 866
rect 838 855 848 858
rect 845 830 848 855
rect 828 826 832 829
rect 841 827 848 830
rect 838 821 841 826
rect 810 818 818 821
rect 793 810 803 813
rect 800 785 803 810
rect 783 781 787 784
rect 796 782 803 785
rect 793 776 796 781
rect 765 773 773 776
rect 748 765 758 768
rect 755 740 758 765
rect 738 736 742 739
rect 751 737 758 740
rect 748 731 751 736
rect 720 728 728 731
rect 703 720 713 723
rect 710 695 713 720
rect 693 691 697 694
rect 706 692 713 695
rect 703 686 706 691
rect 675 683 683 686
rect 658 675 668 678
rect 665 650 668 675
rect 648 646 652 649
rect 661 647 668 650
rect 658 641 661 646
rect 630 638 638 641
rect 613 630 623 633
rect 620 605 623 630
rect 603 601 607 604
rect 616 602 623 605
rect 613 596 616 601
rect 585 593 593 596
rect 568 585 578 588
rect 575 560 578 585
rect 558 556 562 559
rect 571 557 578 560
rect 568 551 571 556
rect 540 548 548 551
rect 523 540 533 543
rect 530 515 533 540
rect 513 511 517 514
rect 526 512 533 515
rect 523 506 526 511
rect 495 503 503 506
rect 478 495 488 498
rect 485 470 488 495
rect 468 466 472 469
rect 481 467 488 470
rect 478 461 481 466
rect 450 458 458 461
rect 433 450 443 453
rect 440 425 443 450
rect 423 421 427 424
rect 436 422 443 425
rect 433 416 436 421
rect 405 413 413 416
rect 388 405 398 408
rect 395 380 398 405
rect 378 376 382 379
rect 391 377 398 380
rect 388 371 391 376
rect 360 368 368 371
rect 343 360 353 363
rect 350 335 353 360
rect 333 331 337 334
rect 346 332 353 335
rect 343 326 346 331
rect 315 323 323 326
rect 298 315 308 318
rect 305 290 308 315
rect 288 286 292 289
rect 301 287 308 290
rect 298 281 301 286
rect 270 278 278 281
rect 253 270 263 273
rect 260 245 263 270
rect 243 241 247 244
rect 256 242 263 245
rect 253 236 256 241
rect 225 233 233 236
rect 208 225 218 228
rect 215 200 218 225
rect 198 196 202 199
rect 211 197 218 200
rect 208 191 211 196
rect 180 188 188 191
rect 163 180 173 183
rect 170 155 173 180
rect 153 151 157 154
rect 166 152 173 155
rect 163 146 166 151
rect 135 143 143 146
rect 118 135 128 138
rect 125 110 128 135
rect 108 106 112 109
rect 121 107 128 110
rect 118 101 121 106
rect 90 98 98 101
rect 73 90 83 93
rect 80 65 83 90
rect 63 61 67 64
rect 76 62 83 65
rect 73 56 76 61
rect 45 53 53 56
rect 28 45 38 48
rect 35 20 38 45
rect 18 16 22 19
rect 31 17 38 20
rect 28 11 31 16
rect 0 8 8 11
rect 0 0 3 8
rect 28 3 31 7
rect 45 11 48 53
rect 73 48 76 52
rect 90 56 93 98
rect 118 93 121 97
rect 135 101 138 143
rect 163 138 166 142
rect 180 146 183 188
rect 208 183 211 187
rect 225 191 228 233
rect 253 228 256 232
rect 270 236 273 278
rect 298 273 301 277
rect 315 281 318 323
rect 343 318 346 322
rect 360 326 363 368
rect 388 363 391 367
rect 405 371 408 413
rect 433 408 436 412
rect 450 416 453 458
rect 478 453 481 457
rect 495 461 498 503
rect 523 498 526 502
rect 540 506 543 548
rect 568 543 571 547
rect 585 551 588 593
rect 613 588 616 592
rect 630 596 633 638
rect 658 633 661 637
rect 675 641 678 683
rect 703 678 706 682
rect 720 686 723 728
rect 748 723 751 727
rect 765 731 768 773
rect 793 768 796 772
rect 810 776 813 818
rect 838 813 841 817
rect 855 821 858 863
rect 883 858 886 862
rect 883 855 893 858
rect 890 830 893 855
rect 873 826 877 829
rect 886 827 893 830
rect 883 821 886 826
rect 855 818 863 821
rect 838 810 848 813
rect 845 785 848 810
rect 828 781 832 784
rect 841 782 848 785
rect 838 776 841 781
rect 810 773 818 776
rect 793 765 803 768
rect 800 740 803 765
rect 783 736 787 739
rect 796 737 803 740
rect 793 731 796 736
rect 765 728 773 731
rect 748 720 758 723
rect 755 695 758 720
rect 738 691 742 694
rect 751 692 758 695
rect 748 686 751 691
rect 720 683 728 686
rect 703 675 713 678
rect 710 650 713 675
rect 693 646 697 649
rect 706 647 713 650
rect 703 641 706 646
rect 675 638 683 641
rect 658 630 668 633
rect 665 605 668 630
rect 648 601 652 604
rect 661 602 668 605
rect 658 596 661 601
rect 630 593 638 596
rect 613 585 623 588
rect 620 560 623 585
rect 603 556 607 559
rect 616 557 623 560
rect 613 551 616 556
rect 585 548 593 551
rect 568 540 578 543
rect 575 515 578 540
rect 558 511 562 514
rect 571 512 578 515
rect 568 506 571 511
rect 540 503 548 506
rect 523 495 533 498
rect 530 470 533 495
rect 513 466 517 469
rect 526 467 533 470
rect 523 461 526 466
rect 495 458 503 461
rect 478 450 488 453
rect 485 425 488 450
rect 468 421 472 424
rect 481 422 488 425
rect 478 416 481 421
rect 450 413 458 416
rect 433 405 443 408
rect 440 380 443 405
rect 423 376 427 379
rect 436 377 443 380
rect 433 371 436 376
rect 405 368 413 371
rect 388 360 398 363
rect 395 335 398 360
rect 378 331 382 334
rect 391 332 398 335
rect 388 326 391 331
rect 360 323 368 326
rect 343 315 353 318
rect 350 290 353 315
rect 333 286 337 289
rect 346 287 353 290
rect 343 281 346 286
rect 315 278 323 281
rect 298 270 308 273
rect 305 245 308 270
rect 288 241 292 244
rect 301 242 308 245
rect 298 236 301 241
rect 270 233 278 236
rect 253 225 263 228
rect 260 200 263 225
rect 243 196 247 199
rect 256 197 263 200
rect 253 191 256 196
rect 225 188 233 191
rect 208 180 218 183
rect 215 155 218 180
rect 198 151 202 154
rect 211 152 218 155
rect 208 146 211 151
rect 180 143 188 146
rect 163 135 173 138
rect 170 110 173 135
rect 153 106 157 109
rect 166 107 173 110
rect 163 101 166 106
rect 135 98 143 101
rect 118 90 128 93
rect 125 65 128 90
rect 108 61 112 64
rect 121 62 128 65
rect 118 56 121 61
rect 90 53 98 56
rect 73 45 83 48
rect 80 20 83 45
rect 63 16 67 19
rect 76 17 83 20
rect 73 11 76 16
rect 45 8 53 11
rect 28 0 38 3
rect 45 0 48 8
rect 73 3 76 7
rect 90 11 93 53
rect 118 48 121 52
rect 135 56 138 98
rect 163 93 166 97
rect 180 101 183 143
rect 208 138 211 142
rect 225 146 228 188
rect 253 183 256 187
rect 270 191 273 233
rect 298 228 301 232
rect 315 236 318 278
rect 343 273 346 277
rect 360 281 363 323
rect 388 318 391 322
rect 405 326 408 368
rect 433 363 436 367
rect 450 371 453 413
rect 478 408 481 412
rect 495 416 498 458
rect 523 453 526 457
rect 540 461 543 503
rect 568 498 571 502
rect 585 506 588 548
rect 613 543 616 547
rect 630 551 633 593
rect 658 588 661 592
rect 675 596 678 638
rect 703 633 706 637
rect 720 641 723 683
rect 748 678 751 682
rect 765 686 768 728
rect 793 723 796 727
rect 810 731 813 773
rect 838 768 841 772
rect 855 776 858 818
rect 883 813 886 817
rect 883 810 893 813
rect 890 785 893 810
rect 873 781 877 784
rect 886 782 893 785
rect 883 776 886 781
rect 855 773 863 776
rect 838 765 848 768
rect 845 740 848 765
rect 828 736 832 739
rect 841 737 848 740
rect 838 731 841 736
rect 810 728 818 731
rect 793 720 803 723
rect 800 695 803 720
rect 783 691 787 694
rect 796 692 803 695
rect 793 686 796 691
rect 765 683 773 686
rect 748 675 758 678
rect 755 650 758 675
rect 738 646 742 649
rect 751 647 758 650
rect 748 641 751 646
rect 720 638 728 641
rect 703 630 713 633
rect 710 605 713 630
rect 693 601 697 604
rect 706 602 713 605
rect 703 596 706 601
rect 675 593 683 596
rect 658 585 668 588
rect 665 560 668 585
rect 648 556 652 559
rect 661 557 668 560
rect 658 551 661 556
rect 630 548 638 551
rect 613 540 623 543
rect 620 515 623 540
rect 603 511 607 514
rect 616 512 623 515
rect 613 506 616 511
rect 585 503 593 506
rect 568 495 578 498
rect 575 470 578 495
rect 558 466 562 469
rect 571 467 578 470
rect 568 461 571 466
rect 540 458 548 461
rect 523 450 533 453
rect 530 425 533 450
rect 513 421 517 424
rect 526 422 533 425
rect 523 416 526 421
rect 495 413 503 416
rect 478 405 488 408
rect 485 380 488 405
rect 468 376 472 379
rect 481 377 488 380
rect 478 371 481 376
rect 450 368 458 371
rect 433 360 443 363
rect 440 335 443 360
rect 423 331 427 334
rect 436 332 443 335
rect 433 326 436 331
rect 405 323 413 326
rect 388 315 398 318
rect 395 290 398 315
rect 378 286 382 289
rect 391 287 398 290
rect 388 281 391 286
rect 360 278 368 281
rect 343 270 353 273
rect 350 245 353 270
rect 333 241 337 244
rect 346 242 353 245
rect 343 236 346 241
rect 315 233 323 236
rect 298 225 308 228
rect 305 200 308 225
rect 288 196 292 199
rect 301 197 308 200
rect 298 191 301 196
rect 270 188 278 191
rect 253 180 263 183
rect 260 155 263 180
rect 243 151 247 154
rect 256 152 263 155
rect 253 146 256 151
rect 225 143 233 146
rect 208 135 218 138
rect 215 110 218 135
rect 198 106 202 109
rect 211 107 218 110
rect 208 101 211 106
rect 180 98 188 101
rect 163 90 173 93
rect 170 65 173 90
rect 153 61 157 64
rect 166 62 173 65
rect 163 56 166 61
rect 135 53 143 56
rect 118 45 128 48
rect 125 20 128 45
rect 108 16 112 19
rect 121 17 128 20
rect 118 11 121 16
rect 90 8 98 11
rect 73 0 83 3
rect 90 0 93 8
rect 118 3 121 7
rect 135 11 138 53
rect 163 48 166 52
rect 180 56 183 98
rect 208 93 211 97
rect 225 101 228 143
rect 253 138 256 142
rect 270 146 273 188
rect 298 183 301 187
rect 315 191 318 233
rect 343 228 346 232
rect 360 236 363 278
rect 388 273 391 277
rect 405 281 408 323
rect 433 318 436 322
rect 450 326 453 368
rect 478 363 481 367
rect 495 371 498 413
rect 523 408 526 412
rect 540 416 543 458
rect 568 453 571 457
rect 585 461 588 503
rect 613 498 616 502
rect 630 506 633 548
rect 658 543 661 547
rect 675 551 678 593
rect 703 588 706 592
rect 720 596 723 638
rect 748 633 751 637
rect 765 641 768 683
rect 793 678 796 682
rect 810 686 813 728
rect 838 723 841 727
rect 855 731 858 773
rect 883 768 886 772
rect 883 765 893 768
rect 890 740 893 765
rect 873 736 877 739
rect 886 737 893 740
rect 883 731 886 736
rect 855 728 863 731
rect 838 720 848 723
rect 845 695 848 720
rect 828 691 832 694
rect 841 692 848 695
rect 838 686 841 691
rect 810 683 818 686
rect 793 675 803 678
rect 800 650 803 675
rect 783 646 787 649
rect 796 647 803 650
rect 793 641 796 646
rect 765 638 773 641
rect 748 630 758 633
rect 755 605 758 630
rect 738 601 742 604
rect 751 602 758 605
rect 748 596 751 601
rect 720 593 728 596
rect 703 585 713 588
rect 710 560 713 585
rect 693 556 697 559
rect 706 557 713 560
rect 703 551 706 556
rect 675 548 683 551
rect 658 540 668 543
rect 665 515 668 540
rect 648 511 652 514
rect 661 512 668 515
rect 658 506 661 511
rect 630 503 638 506
rect 613 495 623 498
rect 620 470 623 495
rect 603 466 607 469
rect 616 467 623 470
rect 613 461 616 466
rect 585 458 593 461
rect 568 450 578 453
rect 575 425 578 450
rect 558 421 562 424
rect 571 422 578 425
rect 568 416 571 421
rect 540 413 548 416
rect 523 405 533 408
rect 530 380 533 405
rect 513 376 517 379
rect 526 377 533 380
rect 523 371 526 376
rect 495 368 503 371
rect 478 360 488 363
rect 485 335 488 360
rect 468 331 472 334
rect 481 332 488 335
rect 478 326 481 331
rect 450 323 458 326
rect 433 315 443 318
rect 440 290 443 315
rect 423 286 427 289
rect 436 287 443 290
rect 433 281 436 286
rect 405 278 413 281
rect 388 270 398 273
rect 395 245 398 270
rect 378 241 382 244
rect 391 242 398 245
rect 388 236 391 241
rect 360 233 368 236
rect 343 225 353 228
rect 350 200 353 225
rect 333 196 337 199
rect 346 197 353 200
rect 343 191 346 196
rect 315 188 323 191
rect 298 180 308 183
rect 305 155 308 180
rect 288 151 292 154
rect 301 152 308 155
rect 298 146 301 151
rect 270 143 278 146
rect 253 135 263 138
rect 260 110 263 135
rect 243 106 247 109
rect 256 107 263 110
rect 253 101 256 106
rect 225 98 233 101
rect 208 90 218 93
rect 215 65 218 90
rect 198 61 202 64
rect 211 62 218 65
rect 208 56 211 61
rect 180 53 188 56
rect 163 45 173 48
rect 170 20 173 45
rect 153 16 157 19
rect 166 17 173 20
rect 163 11 166 16
rect 135 8 143 11
rect 118 0 128 3
rect 135 0 138 8
rect 163 3 166 7
rect 180 11 183 53
rect 208 48 211 52
rect 225 56 228 98
rect 253 93 256 97
rect 270 101 273 143
rect 298 138 301 142
rect 315 146 318 188
rect 343 183 346 187
rect 360 191 363 233
rect 388 228 391 232
rect 405 236 408 278
rect 433 273 436 277
rect 450 281 453 323
rect 478 318 481 322
rect 495 326 498 368
rect 523 363 526 367
rect 540 371 543 413
rect 568 408 571 412
rect 585 416 588 458
rect 613 453 616 457
rect 630 461 633 503
rect 658 498 661 502
rect 675 506 678 548
rect 703 543 706 547
rect 720 551 723 593
rect 748 588 751 592
rect 765 596 768 638
rect 793 633 796 637
rect 810 641 813 683
rect 838 678 841 682
rect 855 686 858 728
rect 883 723 886 727
rect 883 720 893 723
rect 890 695 893 720
rect 873 691 877 694
rect 886 692 893 695
rect 883 686 886 691
rect 855 683 863 686
rect 838 675 848 678
rect 845 650 848 675
rect 828 646 832 649
rect 841 647 848 650
rect 838 641 841 646
rect 810 638 818 641
rect 793 630 803 633
rect 800 605 803 630
rect 783 601 787 604
rect 796 602 803 605
rect 793 596 796 601
rect 765 593 773 596
rect 748 585 758 588
rect 755 560 758 585
rect 738 556 742 559
rect 751 557 758 560
rect 748 551 751 556
rect 720 548 728 551
rect 703 540 713 543
rect 710 515 713 540
rect 693 511 697 514
rect 706 512 713 515
rect 703 506 706 511
rect 675 503 683 506
rect 658 495 668 498
rect 665 470 668 495
rect 648 466 652 469
rect 661 467 668 470
rect 658 461 661 466
rect 630 458 638 461
rect 613 450 623 453
rect 620 425 623 450
rect 603 421 607 424
rect 616 422 623 425
rect 613 416 616 421
rect 585 413 593 416
rect 568 405 578 408
rect 575 380 578 405
rect 558 376 562 379
rect 571 377 578 380
rect 568 371 571 376
rect 540 368 548 371
rect 523 360 533 363
rect 530 335 533 360
rect 513 331 517 334
rect 526 332 533 335
rect 523 326 526 331
rect 495 323 503 326
rect 478 315 488 318
rect 485 290 488 315
rect 468 286 472 289
rect 481 287 488 290
rect 478 281 481 286
rect 450 278 458 281
rect 433 270 443 273
rect 440 245 443 270
rect 423 241 427 244
rect 436 242 443 245
rect 433 236 436 241
rect 405 233 413 236
rect 388 225 398 228
rect 395 200 398 225
rect 378 196 382 199
rect 391 197 398 200
rect 388 191 391 196
rect 360 188 368 191
rect 343 180 353 183
rect 350 155 353 180
rect 333 151 337 154
rect 346 152 353 155
rect 343 146 346 151
rect 315 143 323 146
rect 298 135 308 138
rect 305 110 308 135
rect 288 106 292 109
rect 301 107 308 110
rect 298 101 301 106
rect 270 98 278 101
rect 253 90 263 93
rect 260 65 263 90
rect 243 61 247 64
rect 256 62 263 65
rect 253 56 256 61
rect 225 53 233 56
rect 208 45 218 48
rect 215 20 218 45
rect 198 16 202 19
rect 211 17 218 20
rect 208 11 211 16
rect 180 8 188 11
rect 163 0 173 3
rect 180 0 183 8
rect 208 3 211 7
rect 225 11 228 53
rect 253 48 256 52
rect 270 56 273 98
rect 298 93 301 97
rect 315 101 318 143
rect 343 138 346 142
rect 360 146 363 188
rect 388 183 391 187
rect 405 191 408 233
rect 433 228 436 232
rect 450 236 453 278
rect 478 273 481 277
rect 495 281 498 323
rect 523 318 526 322
rect 540 326 543 368
rect 568 363 571 367
rect 585 371 588 413
rect 613 408 616 412
rect 630 416 633 458
rect 658 453 661 457
rect 675 461 678 503
rect 703 498 706 502
rect 720 506 723 548
rect 748 543 751 547
rect 765 551 768 593
rect 793 588 796 592
rect 810 596 813 638
rect 838 633 841 637
rect 855 641 858 683
rect 883 678 886 682
rect 883 675 893 678
rect 890 650 893 675
rect 873 646 877 649
rect 886 647 893 650
rect 883 641 886 646
rect 855 638 863 641
rect 838 630 848 633
rect 845 605 848 630
rect 828 601 832 604
rect 841 602 848 605
rect 838 596 841 601
rect 810 593 818 596
rect 793 585 803 588
rect 800 560 803 585
rect 783 556 787 559
rect 796 557 803 560
rect 793 551 796 556
rect 765 548 773 551
rect 748 540 758 543
rect 755 515 758 540
rect 738 511 742 514
rect 751 512 758 515
rect 748 506 751 511
rect 720 503 728 506
rect 703 495 713 498
rect 710 470 713 495
rect 693 466 697 469
rect 706 467 713 470
rect 703 461 706 466
rect 675 458 683 461
rect 658 450 668 453
rect 665 425 668 450
rect 648 421 652 424
rect 661 422 668 425
rect 658 416 661 421
rect 630 413 638 416
rect 613 405 623 408
rect 620 380 623 405
rect 603 376 607 379
rect 616 377 623 380
rect 613 371 616 376
rect 585 368 593 371
rect 568 360 578 363
rect 575 335 578 360
rect 558 331 562 334
rect 571 332 578 335
rect 568 326 571 331
rect 540 323 548 326
rect 523 315 533 318
rect 530 290 533 315
rect 513 286 517 289
rect 526 287 533 290
rect 523 281 526 286
rect 495 278 503 281
rect 478 270 488 273
rect 485 245 488 270
rect 468 241 472 244
rect 481 242 488 245
rect 478 236 481 241
rect 450 233 458 236
rect 433 225 443 228
rect 440 200 443 225
rect 423 196 427 199
rect 436 197 443 200
rect 433 191 436 196
rect 405 188 413 191
rect 388 180 398 183
rect 395 155 398 180
rect 378 151 382 154
rect 391 152 398 155
rect 388 146 391 151
rect 360 143 368 146
rect 343 135 353 138
rect 350 110 353 135
rect 333 106 337 109
rect 346 107 353 110
rect 343 101 346 106
rect 315 98 323 101
rect 298 90 308 93
rect 305 65 308 90
rect 288 61 292 64
rect 301 62 308 65
rect 298 56 301 61
rect 270 53 278 56
rect 253 45 263 48
rect 260 20 263 45
rect 243 16 247 19
rect 256 17 263 20
rect 253 11 256 16
rect 225 8 233 11
rect 208 0 218 3
rect 225 0 228 8
rect 253 3 256 7
rect 270 11 273 53
rect 298 48 301 52
rect 315 56 318 98
rect 343 93 346 97
rect 360 101 363 143
rect 388 138 391 142
rect 405 146 408 188
rect 433 183 436 187
rect 450 191 453 233
rect 478 228 481 232
rect 495 236 498 278
rect 523 273 526 277
rect 540 281 543 323
rect 568 318 571 322
rect 585 326 588 368
rect 613 363 616 367
rect 630 371 633 413
rect 658 408 661 412
rect 675 416 678 458
rect 703 453 706 457
rect 720 461 723 503
rect 748 498 751 502
rect 765 506 768 548
rect 793 543 796 547
rect 810 551 813 593
rect 838 588 841 592
rect 855 596 858 638
rect 883 633 886 637
rect 883 630 893 633
rect 890 605 893 630
rect 873 601 877 604
rect 886 602 893 605
rect 883 596 886 601
rect 855 593 863 596
rect 838 585 848 588
rect 845 560 848 585
rect 828 556 832 559
rect 841 557 848 560
rect 838 551 841 556
rect 810 548 818 551
rect 793 540 803 543
rect 800 515 803 540
rect 783 511 787 514
rect 796 512 803 515
rect 793 506 796 511
rect 765 503 773 506
rect 748 495 758 498
rect 755 470 758 495
rect 738 466 742 469
rect 751 467 758 470
rect 748 461 751 466
rect 720 458 728 461
rect 703 450 713 453
rect 710 425 713 450
rect 693 421 697 424
rect 706 422 713 425
rect 703 416 706 421
rect 675 413 683 416
rect 658 405 668 408
rect 665 380 668 405
rect 648 376 652 379
rect 661 377 668 380
rect 658 371 661 376
rect 630 368 638 371
rect 613 360 623 363
rect 620 335 623 360
rect 603 331 607 334
rect 616 332 623 335
rect 613 326 616 331
rect 585 323 593 326
rect 568 315 578 318
rect 575 290 578 315
rect 558 286 562 289
rect 571 287 578 290
rect 568 281 571 286
rect 540 278 548 281
rect 523 270 533 273
rect 530 245 533 270
rect 513 241 517 244
rect 526 242 533 245
rect 523 236 526 241
rect 495 233 503 236
rect 478 225 488 228
rect 485 200 488 225
rect 468 196 472 199
rect 481 197 488 200
rect 478 191 481 196
rect 450 188 458 191
rect 433 180 443 183
rect 440 155 443 180
rect 423 151 427 154
rect 436 152 443 155
rect 433 146 436 151
rect 405 143 413 146
rect 388 135 398 138
rect 395 110 398 135
rect 378 106 382 109
rect 391 107 398 110
rect 388 101 391 106
rect 360 98 368 101
rect 343 90 353 93
rect 350 65 353 90
rect 333 61 337 64
rect 346 62 353 65
rect 343 56 346 61
rect 315 53 323 56
rect 298 45 308 48
rect 305 20 308 45
rect 288 16 292 19
rect 301 17 308 20
rect 298 11 301 16
rect 270 8 278 11
rect 253 0 263 3
rect 270 0 273 8
rect 298 3 301 7
rect 315 11 318 53
rect 343 48 346 52
rect 360 56 363 98
rect 388 93 391 97
rect 405 101 408 143
rect 433 138 436 142
rect 450 146 453 188
rect 478 183 481 187
rect 495 191 498 233
rect 523 228 526 232
rect 540 236 543 278
rect 568 273 571 277
rect 585 281 588 323
rect 613 318 616 322
rect 630 326 633 368
rect 658 363 661 367
rect 675 371 678 413
rect 703 408 706 412
rect 720 416 723 458
rect 748 453 751 457
rect 765 461 768 503
rect 793 498 796 502
rect 810 506 813 548
rect 838 543 841 547
rect 855 551 858 593
rect 883 588 886 592
rect 883 585 893 588
rect 890 560 893 585
rect 873 556 877 559
rect 886 557 893 560
rect 883 551 886 556
rect 855 548 863 551
rect 838 540 848 543
rect 845 515 848 540
rect 828 511 832 514
rect 841 512 848 515
rect 838 506 841 511
rect 810 503 818 506
rect 793 495 803 498
rect 800 470 803 495
rect 783 466 787 469
rect 796 467 803 470
rect 793 461 796 466
rect 765 458 773 461
rect 748 450 758 453
rect 755 425 758 450
rect 738 421 742 424
rect 751 422 758 425
rect 748 416 751 421
rect 720 413 728 416
rect 703 405 713 408
rect 710 380 713 405
rect 693 376 697 379
rect 706 377 713 380
rect 703 371 706 376
rect 675 368 683 371
rect 658 360 668 363
rect 665 335 668 360
rect 648 331 652 334
rect 661 332 668 335
rect 658 326 661 331
rect 630 323 638 326
rect 613 315 623 318
rect 620 290 623 315
rect 603 286 607 289
rect 616 287 623 290
rect 613 281 616 286
rect 585 278 593 281
rect 568 270 578 273
rect 575 245 578 270
rect 558 241 562 244
rect 571 242 578 245
rect 568 236 571 241
rect 540 233 548 236
rect 523 225 533 228
rect 530 200 533 225
rect 513 196 517 199
rect 526 197 533 200
rect 523 191 526 196
rect 495 188 503 191
rect 478 180 488 183
rect 485 155 488 180
rect 468 151 472 154
rect 481 152 488 155
rect 478 146 481 151
rect 450 143 458 146
rect 433 135 443 138
rect 440 110 443 135
rect 423 106 427 109
rect 436 107 443 110
rect 433 101 436 106
rect 405 98 413 101
rect 388 90 398 93
rect 395 65 398 90
rect 378 61 382 64
rect 391 62 398 65
rect 388 56 391 61
rect 360 53 368 56
rect 343 45 353 48
rect 350 20 353 45
rect 333 16 337 19
rect 346 17 353 20
rect 343 11 346 16
rect 315 8 323 11
rect 298 0 308 3
rect 315 0 318 8
rect 343 3 346 7
rect 360 11 363 53
rect 388 48 391 52
rect 405 56 408 98
rect 433 93 436 97
rect 450 101 453 143
rect 478 138 481 142
rect 495 146 498 188
rect 523 183 526 187
rect 540 191 543 233
rect 568 228 571 232
rect 585 236 588 278
rect 613 273 616 277
rect 630 281 633 323
rect 658 318 661 322
rect 675 326 678 368
rect 703 363 706 367
rect 720 371 723 413
rect 748 408 751 412
rect 765 416 768 458
rect 793 453 796 457
rect 810 461 813 503
rect 838 498 841 502
rect 855 506 858 548
rect 883 543 886 547
rect 883 540 893 543
rect 890 515 893 540
rect 873 511 877 514
rect 886 512 893 515
rect 883 506 886 511
rect 855 503 863 506
rect 838 495 848 498
rect 845 470 848 495
rect 828 466 832 469
rect 841 467 848 470
rect 838 461 841 466
rect 810 458 818 461
rect 793 450 803 453
rect 800 425 803 450
rect 783 421 787 424
rect 796 422 803 425
rect 793 416 796 421
rect 765 413 773 416
rect 748 405 758 408
rect 755 380 758 405
rect 738 376 742 379
rect 751 377 758 380
rect 748 371 751 376
rect 720 368 728 371
rect 703 360 713 363
rect 710 335 713 360
rect 693 331 697 334
rect 706 332 713 335
rect 703 326 706 331
rect 675 323 683 326
rect 658 315 668 318
rect 665 290 668 315
rect 648 286 652 289
rect 661 287 668 290
rect 658 281 661 286
rect 630 278 638 281
rect 613 270 623 273
rect 620 245 623 270
rect 603 241 607 244
rect 616 242 623 245
rect 613 236 616 241
rect 585 233 593 236
rect 568 225 578 228
rect 575 200 578 225
rect 558 196 562 199
rect 571 197 578 200
rect 568 191 571 196
rect 540 188 548 191
rect 523 180 533 183
rect 530 155 533 180
rect 513 151 517 154
rect 526 152 533 155
rect 523 146 526 151
rect 495 143 503 146
rect 478 135 488 138
rect 485 110 488 135
rect 468 106 472 109
rect 481 107 488 110
rect 478 101 481 106
rect 450 98 458 101
rect 433 90 443 93
rect 440 65 443 90
rect 423 61 427 64
rect 436 62 443 65
rect 433 56 436 61
rect 405 53 413 56
rect 388 45 398 48
rect 395 20 398 45
rect 378 16 382 19
rect 391 17 398 20
rect 388 11 391 16
rect 360 8 368 11
rect 343 0 353 3
rect 360 0 363 8
rect 388 3 391 7
rect 405 11 408 53
rect 433 48 436 52
rect 450 56 453 98
rect 478 93 481 97
rect 495 101 498 143
rect 523 138 526 142
rect 540 146 543 188
rect 568 183 571 187
rect 585 191 588 233
rect 613 228 616 232
rect 630 236 633 278
rect 658 273 661 277
rect 675 281 678 323
rect 703 318 706 322
rect 720 326 723 368
rect 748 363 751 367
rect 765 371 768 413
rect 793 408 796 412
rect 810 416 813 458
rect 838 453 841 457
rect 855 461 858 503
rect 883 498 886 502
rect 883 495 893 498
rect 890 470 893 495
rect 873 466 877 469
rect 886 467 893 470
rect 883 461 886 466
rect 855 458 863 461
rect 838 450 848 453
rect 845 425 848 450
rect 828 421 832 424
rect 841 422 848 425
rect 838 416 841 421
rect 810 413 818 416
rect 793 405 803 408
rect 800 380 803 405
rect 783 376 787 379
rect 796 377 803 380
rect 793 371 796 376
rect 765 368 773 371
rect 748 360 758 363
rect 755 335 758 360
rect 738 331 742 334
rect 751 332 758 335
rect 748 326 751 331
rect 720 323 728 326
rect 703 315 713 318
rect 710 290 713 315
rect 693 286 697 289
rect 706 287 713 290
rect 703 281 706 286
rect 675 278 683 281
rect 658 270 668 273
rect 665 245 668 270
rect 648 241 652 244
rect 661 242 668 245
rect 658 236 661 241
rect 630 233 638 236
rect 613 225 623 228
rect 620 200 623 225
rect 603 196 607 199
rect 616 197 623 200
rect 613 191 616 196
rect 585 188 593 191
rect 568 180 578 183
rect 575 155 578 180
rect 558 151 562 154
rect 571 152 578 155
rect 568 146 571 151
rect 540 143 548 146
rect 523 135 533 138
rect 530 110 533 135
rect 513 106 517 109
rect 526 107 533 110
rect 523 101 526 106
rect 495 98 503 101
rect 478 90 488 93
rect 485 65 488 90
rect 468 61 472 64
rect 481 62 488 65
rect 478 56 481 61
rect 450 53 458 56
rect 433 45 443 48
rect 440 20 443 45
rect 423 16 427 19
rect 436 17 443 20
rect 433 11 436 16
rect 405 8 413 11
rect 388 0 398 3
rect 405 0 408 8
rect 433 3 436 7
rect 450 11 453 53
rect 478 48 481 52
rect 495 56 498 98
rect 523 93 526 97
rect 540 101 543 143
rect 568 138 571 142
rect 585 146 588 188
rect 613 183 616 187
rect 630 191 633 233
rect 658 228 661 232
rect 675 236 678 278
rect 703 273 706 277
rect 720 281 723 323
rect 748 318 751 322
rect 765 326 768 368
rect 793 363 796 367
rect 810 371 813 413
rect 838 408 841 412
rect 855 416 858 458
rect 883 453 886 457
rect 883 450 893 453
rect 890 425 893 450
rect 873 421 877 424
rect 886 422 893 425
rect 883 416 886 421
rect 855 413 863 416
rect 838 405 848 408
rect 845 380 848 405
rect 828 376 832 379
rect 841 377 848 380
rect 838 371 841 376
rect 810 368 818 371
rect 793 360 803 363
rect 800 335 803 360
rect 783 331 787 334
rect 796 332 803 335
rect 793 326 796 331
rect 765 323 773 326
rect 748 315 758 318
rect 755 290 758 315
rect 738 286 742 289
rect 751 287 758 290
rect 748 281 751 286
rect 720 278 728 281
rect 703 270 713 273
rect 710 245 713 270
rect 693 241 697 244
rect 706 242 713 245
rect 703 236 706 241
rect 675 233 683 236
rect 658 225 668 228
rect 665 200 668 225
rect 648 196 652 199
rect 661 197 668 200
rect 658 191 661 196
rect 630 188 638 191
rect 613 180 623 183
rect 620 155 623 180
rect 603 151 607 154
rect 616 152 623 155
rect 613 146 616 151
rect 585 143 593 146
rect 568 135 578 138
rect 575 110 578 135
rect 558 106 562 109
rect 571 107 578 110
rect 568 101 571 106
rect 540 98 548 101
rect 523 90 533 93
rect 530 65 533 90
rect 513 61 517 64
rect 526 62 533 65
rect 523 56 526 61
rect 495 53 503 56
rect 478 45 488 48
rect 485 20 488 45
rect 468 16 472 19
rect 481 17 488 20
rect 478 11 481 16
rect 450 8 458 11
rect 433 0 443 3
rect 450 0 453 8
rect 478 3 481 7
rect 495 11 498 53
rect 523 48 526 52
rect 540 56 543 98
rect 568 93 571 97
rect 585 101 588 143
rect 613 138 616 142
rect 630 146 633 188
rect 658 183 661 187
rect 675 191 678 233
rect 703 228 706 232
rect 720 236 723 278
rect 748 273 751 277
rect 765 281 768 323
rect 793 318 796 322
rect 810 326 813 368
rect 838 363 841 367
rect 855 371 858 413
rect 883 408 886 412
rect 883 405 893 408
rect 890 380 893 405
rect 873 376 877 379
rect 886 377 893 380
rect 883 371 886 376
rect 855 368 863 371
rect 838 360 848 363
rect 845 335 848 360
rect 828 331 832 334
rect 841 332 848 335
rect 838 326 841 331
rect 810 323 818 326
rect 793 315 803 318
rect 800 290 803 315
rect 783 286 787 289
rect 796 287 803 290
rect 793 281 796 286
rect 765 278 773 281
rect 748 270 758 273
rect 755 245 758 270
rect 738 241 742 244
rect 751 242 758 245
rect 748 236 751 241
rect 720 233 728 236
rect 703 225 713 228
rect 710 200 713 225
rect 693 196 697 199
rect 706 197 713 200
rect 703 191 706 196
rect 675 188 683 191
rect 658 180 668 183
rect 665 155 668 180
rect 648 151 652 154
rect 661 152 668 155
rect 658 146 661 151
rect 630 143 638 146
rect 613 135 623 138
rect 620 110 623 135
rect 603 106 607 109
rect 616 107 623 110
rect 613 101 616 106
rect 585 98 593 101
rect 568 90 578 93
rect 575 65 578 90
rect 558 61 562 64
rect 571 62 578 65
rect 568 56 571 61
rect 540 53 548 56
rect 523 45 533 48
rect 530 20 533 45
rect 513 16 517 19
rect 526 17 533 20
rect 523 11 526 16
rect 495 8 503 11
rect 478 0 488 3
rect 495 0 498 8
rect 523 3 526 7
rect 540 11 543 53
rect 568 48 571 52
rect 585 56 588 98
rect 613 93 616 97
rect 630 101 633 143
rect 658 138 661 142
rect 675 146 678 188
rect 703 183 706 187
rect 720 191 723 233
rect 748 228 751 232
rect 765 236 768 278
rect 793 273 796 277
rect 810 281 813 323
rect 838 318 841 322
rect 855 326 858 368
rect 883 363 886 367
rect 883 360 893 363
rect 890 335 893 360
rect 873 331 877 334
rect 886 332 893 335
rect 883 326 886 331
rect 855 323 863 326
rect 838 315 848 318
rect 845 290 848 315
rect 828 286 832 289
rect 841 287 848 290
rect 838 281 841 286
rect 810 278 818 281
rect 793 270 803 273
rect 800 245 803 270
rect 783 241 787 244
rect 796 242 803 245
rect 793 236 796 241
rect 765 233 773 236
rect 748 225 758 228
rect 755 200 758 225
rect 738 196 742 199
rect 751 197 758 200
rect 748 191 751 196
rect 720 188 728 191
rect 703 180 713 183
rect 710 155 713 180
rect 693 151 697 154
rect 706 152 713 155
rect 703 146 706 151
rect 675 143 683 146
rect 658 135 668 138
rect 665 110 668 135
rect 648 106 652 109
rect 661 107 668 110
rect 658 101 661 106
rect 630 98 638 101
rect 613 90 623 93
rect 620 65 623 90
rect 603 61 607 64
rect 616 62 623 65
rect 613 56 616 61
rect 585 53 593 56
rect 568 45 578 48
rect 575 20 578 45
rect 558 16 562 19
rect 571 17 578 20
rect 568 11 571 16
rect 540 8 548 11
rect 523 0 533 3
rect 540 0 543 8
rect 568 3 571 7
rect 585 11 588 53
rect 613 48 616 52
rect 630 56 633 98
rect 658 93 661 97
rect 675 101 678 143
rect 703 138 706 142
rect 720 146 723 188
rect 748 183 751 187
rect 765 191 768 233
rect 793 228 796 232
rect 810 236 813 278
rect 838 273 841 277
rect 855 281 858 323
rect 883 318 886 322
rect 883 315 893 318
rect 890 290 893 315
rect 873 286 877 289
rect 886 287 893 290
rect 883 281 886 286
rect 855 278 863 281
rect 838 270 848 273
rect 845 245 848 270
rect 828 241 832 244
rect 841 242 848 245
rect 838 236 841 241
rect 810 233 818 236
rect 793 225 803 228
rect 800 200 803 225
rect 783 196 787 199
rect 796 197 803 200
rect 793 191 796 196
rect 765 188 773 191
rect 748 180 758 183
rect 755 155 758 180
rect 738 151 742 154
rect 751 152 758 155
rect 748 146 751 151
rect 720 143 728 146
rect 703 135 713 138
rect 710 110 713 135
rect 693 106 697 109
rect 706 107 713 110
rect 703 101 706 106
rect 675 98 683 101
rect 658 90 668 93
rect 665 65 668 90
rect 648 61 652 64
rect 661 62 668 65
rect 658 56 661 61
rect 630 53 638 56
rect 613 45 623 48
rect 620 20 623 45
rect 603 16 607 19
rect 616 17 623 20
rect 613 11 616 16
rect 585 8 593 11
rect 568 0 578 3
rect 585 0 588 8
rect 613 3 616 7
rect 630 11 633 53
rect 658 48 661 52
rect 675 56 678 98
rect 703 93 706 97
rect 720 101 723 143
rect 748 138 751 142
rect 765 146 768 188
rect 793 183 796 187
rect 810 191 813 233
rect 838 228 841 232
rect 855 236 858 278
rect 883 273 886 277
rect 883 270 893 273
rect 890 245 893 270
rect 873 241 877 244
rect 886 242 893 245
rect 883 236 886 241
rect 855 233 863 236
rect 838 225 848 228
rect 845 200 848 225
rect 828 196 832 199
rect 841 197 848 200
rect 838 191 841 196
rect 810 188 818 191
rect 793 180 803 183
rect 800 155 803 180
rect 783 151 787 154
rect 796 152 803 155
rect 793 146 796 151
rect 765 143 773 146
rect 748 135 758 138
rect 755 110 758 135
rect 738 106 742 109
rect 751 107 758 110
rect 748 101 751 106
rect 720 98 728 101
rect 703 90 713 93
rect 710 65 713 90
rect 693 61 697 64
rect 706 62 713 65
rect 703 56 706 61
rect 675 53 683 56
rect 658 45 668 48
rect 665 20 668 45
rect 648 16 652 19
rect 661 17 668 20
rect 658 11 661 16
rect 630 8 638 11
rect 613 0 623 3
rect 630 0 633 8
rect 658 3 661 7
rect 675 11 678 53
rect 703 48 706 52
rect 720 56 723 98
rect 748 93 751 97
rect 765 101 768 143
rect 793 138 796 142
rect 810 146 813 188
rect 838 183 841 187
rect 855 191 858 233
rect 883 228 886 232
rect 883 225 893 228
rect 890 200 893 225
rect 873 196 877 199
rect 886 197 893 200
rect 883 191 886 196
rect 855 188 863 191
rect 838 180 848 183
rect 845 155 848 180
rect 828 151 832 154
rect 841 152 848 155
rect 838 146 841 151
rect 810 143 818 146
rect 793 135 803 138
rect 800 110 803 135
rect 783 106 787 109
rect 796 107 803 110
rect 793 101 796 106
rect 765 98 773 101
rect 748 90 758 93
rect 755 65 758 90
rect 738 61 742 64
rect 751 62 758 65
rect 748 56 751 61
rect 720 53 728 56
rect 703 45 713 48
rect 710 20 713 45
rect 693 16 697 19
rect 706 17 713 20
rect 703 11 706 16
rect 675 8 683 11
rect 658 0 668 3
rect 675 0 678 8
rect 703 3 706 7
rect 720 11 723 53
rect 748 48 751 52
rect 765 56 768 98
rect 793 93 796 97
rect 810 101 813 143
rect 838 138 841 142
rect 855 146 858 188
rect 883 183 886 187
rect 883 180 893 183
rect 890 155 893 180
rect 873 151 877 154
rect 886 152 893 155
rect 883 146 886 151
rect 855 143 863 146
rect 838 135 848 138
rect 845 110 848 135
rect 828 106 832 109
rect 841 107 848 110
rect 838 101 841 106
rect 810 98 818 101
rect 793 90 803 93
rect 800 65 803 90
rect 783 61 787 64
rect 796 62 803 65
rect 793 56 796 61
rect 765 53 773 56
rect 748 45 758 48
rect 755 20 758 45
rect 738 16 742 19
rect 751 17 758 20
rect 748 11 751 16
rect 720 8 728 11
rect 703 0 713 3
rect 720 0 723 8
rect 748 3 751 7
rect 765 11 768 53
rect 793 48 796 52
rect 810 56 813 98
rect 838 93 841 97
rect 855 101 858 143
rect 883 138 886 142
rect 883 135 893 138
rect 890 110 893 135
rect 873 106 877 109
rect 886 107 893 110
rect 883 101 886 106
rect 855 98 863 101
rect 838 90 848 93
rect 845 65 848 90
rect 828 61 832 64
rect 841 62 848 65
rect 838 56 841 61
rect 810 53 818 56
rect 793 45 803 48
rect 800 20 803 45
rect 783 16 787 19
rect 796 17 803 20
rect 793 11 796 16
rect 765 8 773 11
rect 748 0 758 3
rect 765 0 768 8
rect 793 3 796 7
rect 810 11 813 53
rect 838 48 841 52
rect 855 56 858 98
rect 883 93 886 97
rect 883 90 893 93
rect 890 65 893 90
rect 873 61 877 64
rect 886 62 893 65
rect 883 56 886 61
rect 855 53 863 56
rect 838 45 848 48
rect 845 20 848 45
rect 828 16 832 19
rect 841 17 848 20
rect 838 11 841 16
rect 810 8 818 11
rect 793 0 803 3
rect 810 0 813 8
rect 838 3 841 7
rect 855 11 858 53
rect 883 48 886 52
rect 883 45 893 48
rect 890 20 893 45
rect 873 16 877 19
rect 886 17 893 20
rect 883 11 886 16
rect 855 8 863 11
rect 838 0 848 3
rect 855 0 858 8
rect 883 3 886 7
rect 883 0 893 3
rect -266 -158 -263 -152
rect -296 -172 -293 -168
rect -266 -180 -263 -162
rect -216 -170 -213 -136
rect -181 -161 -178 -136
rect -198 -165 -194 -162
rect -185 -164 -178 -161
rect -188 -170 -185 -165
rect -216 -173 -208 -170
rect -216 -181 -213 -173
rect -188 -178 -185 -174
rect -188 -181 -178 -178
<< m2contact >>
rect 28 878 32 882
rect 19 855 23 859
rect 34 861 38 865
rect 73 878 77 882
rect 28 833 32 837
rect 19 810 23 814
rect 34 816 38 820
rect 64 855 68 859
rect 79 861 83 865
rect 118 878 122 882
rect 73 833 77 837
rect 28 788 32 792
rect 19 765 23 769
rect 34 771 38 775
rect 64 810 68 814
rect 79 816 83 820
rect 109 855 113 859
rect 124 861 128 865
rect 163 878 167 882
rect 118 833 122 837
rect 73 788 77 792
rect 28 743 32 747
rect 19 720 23 724
rect 34 726 38 730
rect 64 765 68 769
rect 79 771 83 775
rect 109 810 113 814
rect 124 816 128 820
rect 154 855 158 859
rect 169 861 173 865
rect 208 878 212 882
rect 163 833 167 837
rect 118 788 122 792
rect 73 743 77 747
rect 28 698 32 702
rect 19 675 23 679
rect 34 681 38 685
rect 64 720 68 724
rect 79 726 83 730
rect 109 765 113 769
rect 124 771 128 775
rect 154 810 158 814
rect 169 816 173 820
rect 199 855 203 859
rect 214 861 218 865
rect 253 878 257 882
rect 208 833 212 837
rect 163 788 167 792
rect 118 743 122 747
rect 73 698 77 702
rect 28 653 32 657
rect 19 630 23 634
rect 34 636 38 640
rect 64 675 68 679
rect 79 681 83 685
rect 109 720 113 724
rect 124 726 128 730
rect 154 765 158 769
rect 169 771 173 775
rect 199 810 203 814
rect 214 816 218 820
rect 244 855 248 859
rect 259 861 263 865
rect 298 878 302 882
rect 253 833 257 837
rect 208 788 212 792
rect 163 743 167 747
rect 118 698 122 702
rect 73 653 77 657
rect 28 608 32 612
rect 19 585 23 589
rect 34 591 38 595
rect 64 630 68 634
rect 79 636 83 640
rect 109 675 113 679
rect 124 681 128 685
rect 154 720 158 724
rect 169 726 173 730
rect 199 765 203 769
rect 214 771 218 775
rect 244 810 248 814
rect 259 816 263 820
rect 289 855 293 859
rect 304 861 308 865
rect 343 878 347 882
rect 298 833 302 837
rect 253 788 257 792
rect 208 743 212 747
rect 163 698 167 702
rect 118 653 122 657
rect 73 608 77 612
rect 28 563 32 567
rect 19 540 23 544
rect 34 546 38 550
rect 64 585 68 589
rect 79 591 83 595
rect 109 630 113 634
rect 124 636 128 640
rect 154 675 158 679
rect 169 681 173 685
rect 199 720 203 724
rect 214 726 218 730
rect 244 765 248 769
rect 259 771 263 775
rect 289 810 293 814
rect 304 816 308 820
rect 334 855 338 859
rect 349 861 353 865
rect 388 878 392 882
rect 343 833 347 837
rect 298 788 302 792
rect 253 743 257 747
rect 208 698 212 702
rect 163 653 167 657
rect 118 608 122 612
rect 73 563 77 567
rect 28 518 32 522
rect 19 495 23 499
rect 34 501 38 505
rect 64 540 68 544
rect 79 546 83 550
rect 109 585 113 589
rect 124 591 128 595
rect 154 630 158 634
rect 169 636 173 640
rect 199 675 203 679
rect 214 681 218 685
rect 244 720 248 724
rect 259 726 263 730
rect 289 765 293 769
rect 304 771 308 775
rect 334 810 338 814
rect 349 816 353 820
rect 379 855 383 859
rect 394 861 398 865
rect 433 878 437 882
rect 388 833 392 837
rect 343 788 347 792
rect 298 743 302 747
rect 253 698 257 702
rect 208 653 212 657
rect 163 608 167 612
rect 118 563 122 567
rect 73 518 77 522
rect 28 473 32 477
rect 19 450 23 454
rect 34 456 38 460
rect 64 495 68 499
rect 79 501 83 505
rect 109 540 113 544
rect 124 546 128 550
rect 154 585 158 589
rect 169 591 173 595
rect 199 630 203 634
rect 214 636 218 640
rect 244 675 248 679
rect 259 681 263 685
rect 289 720 293 724
rect 304 726 308 730
rect 334 765 338 769
rect 349 771 353 775
rect 379 810 383 814
rect 394 816 398 820
rect 424 855 428 859
rect 439 861 443 865
rect 478 878 482 882
rect 433 833 437 837
rect 388 788 392 792
rect 343 743 347 747
rect 298 698 302 702
rect 253 653 257 657
rect 208 608 212 612
rect 163 563 167 567
rect 118 518 122 522
rect 73 473 77 477
rect 28 428 32 432
rect 19 405 23 409
rect 34 411 38 415
rect 64 450 68 454
rect 79 456 83 460
rect 109 495 113 499
rect 124 501 128 505
rect 154 540 158 544
rect 169 546 173 550
rect 199 585 203 589
rect 214 591 218 595
rect 244 630 248 634
rect 259 636 263 640
rect 289 675 293 679
rect 304 681 308 685
rect 334 720 338 724
rect 349 726 353 730
rect 379 765 383 769
rect 394 771 398 775
rect 424 810 428 814
rect 439 816 443 820
rect 469 855 473 859
rect 484 861 488 865
rect 523 878 527 882
rect 478 833 482 837
rect 433 788 437 792
rect 388 743 392 747
rect 343 698 347 702
rect 298 653 302 657
rect 253 608 257 612
rect 208 563 212 567
rect 163 518 167 522
rect 118 473 122 477
rect 73 428 77 432
rect 28 383 32 387
rect 19 360 23 364
rect 34 366 38 370
rect 64 405 68 409
rect 79 411 83 415
rect 109 450 113 454
rect 124 456 128 460
rect 154 495 158 499
rect 169 501 173 505
rect 199 540 203 544
rect 214 546 218 550
rect 244 585 248 589
rect 259 591 263 595
rect 289 630 293 634
rect 304 636 308 640
rect 334 675 338 679
rect 349 681 353 685
rect 379 720 383 724
rect 394 726 398 730
rect 424 765 428 769
rect 439 771 443 775
rect 469 810 473 814
rect 484 816 488 820
rect 514 855 518 859
rect 529 861 533 865
rect 568 878 572 882
rect 523 833 527 837
rect 478 788 482 792
rect 433 743 437 747
rect 388 698 392 702
rect 343 653 347 657
rect 298 608 302 612
rect 253 563 257 567
rect 208 518 212 522
rect 163 473 167 477
rect 118 428 122 432
rect 73 383 77 387
rect 28 338 32 342
rect 19 315 23 319
rect 34 321 38 325
rect 64 360 68 364
rect 79 366 83 370
rect 109 405 113 409
rect 124 411 128 415
rect 154 450 158 454
rect 169 456 173 460
rect 199 495 203 499
rect 214 501 218 505
rect 244 540 248 544
rect 259 546 263 550
rect 289 585 293 589
rect 304 591 308 595
rect 334 630 338 634
rect 349 636 353 640
rect 379 675 383 679
rect 394 681 398 685
rect 424 720 428 724
rect 439 726 443 730
rect 469 765 473 769
rect 484 771 488 775
rect 514 810 518 814
rect 529 816 533 820
rect 559 855 563 859
rect 574 861 578 865
rect 613 878 617 882
rect 568 833 572 837
rect 523 788 527 792
rect 478 743 482 747
rect 433 698 437 702
rect 388 653 392 657
rect 343 608 347 612
rect 298 563 302 567
rect 253 518 257 522
rect 208 473 212 477
rect 163 428 167 432
rect 118 383 122 387
rect 73 338 77 342
rect 28 293 32 297
rect 19 270 23 274
rect 34 276 38 280
rect 64 315 68 319
rect 79 321 83 325
rect 109 360 113 364
rect 124 366 128 370
rect 154 405 158 409
rect 169 411 173 415
rect 199 450 203 454
rect 214 456 218 460
rect 244 495 248 499
rect 259 501 263 505
rect 289 540 293 544
rect 304 546 308 550
rect 334 585 338 589
rect 349 591 353 595
rect 379 630 383 634
rect 394 636 398 640
rect 424 675 428 679
rect 439 681 443 685
rect 469 720 473 724
rect 484 726 488 730
rect 514 765 518 769
rect 529 771 533 775
rect 559 810 563 814
rect 574 816 578 820
rect 604 855 608 859
rect 619 861 623 865
rect 658 878 662 882
rect 613 833 617 837
rect 568 788 572 792
rect 523 743 527 747
rect 478 698 482 702
rect 433 653 437 657
rect 388 608 392 612
rect 343 563 347 567
rect 298 518 302 522
rect 253 473 257 477
rect 208 428 212 432
rect 163 383 167 387
rect 118 338 122 342
rect 73 293 77 297
rect 28 248 32 252
rect 19 225 23 229
rect 34 231 38 235
rect 64 270 68 274
rect 79 276 83 280
rect 109 315 113 319
rect 124 321 128 325
rect 154 360 158 364
rect 169 366 173 370
rect 199 405 203 409
rect 214 411 218 415
rect 244 450 248 454
rect 259 456 263 460
rect 289 495 293 499
rect 304 501 308 505
rect 334 540 338 544
rect 349 546 353 550
rect 379 585 383 589
rect 394 591 398 595
rect 424 630 428 634
rect 439 636 443 640
rect 469 675 473 679
rect 484 681 488 685
rect 514 720 518 724
rect 529 726 533 730
rect 559 765 563 769
rect 574 771 578 775
rect 604 810 608 814
rect 619 816 623 820
rect 649 855 653 859
rect 664 861 668 865
rect 703 878 707 882
rect 658 833 662 837
rect 613 788 617 792
rect 568 743 572 747
rect 523 698 527 702
rect 478 653 482 657
rect 433 608 437 612
rect 388 563 392 567
rect 343 518 347 522
rect 298 473 302 477
rect 253 428 257 432
rect 208 383 212 387
rect 163 338 167 342
rect 118 293 122 297
rect 73 248 77 252
rect 28 203 32 207
rect 19 180 23 184
rect 34 186 38 190
rect 64 225 68 229
rect 79 231 83 235
rect 109 270 113 274
rect 124 276 128 280
rect 154 315 158 319
rect 169 321 173 325
rect 199 360 203 364
rect 214 366 218 370
rect 244 405 248 409
rect 259 411 263 415
rect 289 450 293 454
rect 304 456 308 460
rect 334 495 338 499
rect 349 501 353 505
rect 379 540 383 544
rect 394 546 398 550
rect 424 585 428 589
rect 439 591 443 595
rect 469 630 473 634
rect 484 636 488 640
rect 514 675 518 679
rect 529 681 533 685
rect 559 720 563 724
rect 574 726 578 730
rect 604 765 608 769
rect 619 771 623 775
rect 649 810 653 814
rect 664 816 668 820
rect 694 855 698 859
rect 709 861 713 865
rect 748 878 752 882
rect 703 833 707 837
rect 658 788 662 792
rect 613 743 617 747
rect 568 698 572 702
rect 523 653 527 657
rect 478 608 482 612
rect 433 563 437 567
rect 388 518 392 522
rect 343 473 347 477
rect 298 428 302 432
rect 253 383 257 387
rect 208 338 212 342
rect 163 293 167 297
rect 118 248 122 252
rect 73 203 77 207
rect 28 158 32 162
rect 19 135 23 139
rect 34 141 38 145
rect 64 180 68 184
rect 79 186 83 190
rect 109 225 113 229
rect 124 231 128 235
rect 154 270 158 274
rect 169 276 173 280
rect 199 315 203 319
rect 214 321 218 325
rect 244 360 248 364
rect 259 366 263 370
rect 289 405 293 409
rect 304 411 308 415
rect 334 450 338 454
rect 349 456 353 460
rect 379 495 383 499
rect 394 501 398 505
rect 424 540 428 544
rect 439 546 443 550
rect 469 585 473 589
rect 484 591 488 595
rect 514 630 518 634
rect 529 636 533 640
rect 559 675 563 679
rect 574 681 578 685
rect 604 720 608 724
rect 619 726 623 730
rect 649 765 653 769
rect 664 771 668 775
rect 694 810 698 814
rect 709 816 713 820
rect 739 855 743 859
rect 754 861 758 865
rect 793 878 797 882
rect 748 833 752 837
rect 703 788 707 792
rect 658 743 662 747
rect 613 698 617 702
rect 568 653 572 657
rect 523 608 527 612
rect 478 563 482 567
rect 433 518 437 522
rect 388 473 392 477
rect 343 428 347 432
rect 298 383 302 387
rect 253 338 257 342
rect 208 293 212 297
rect 163 248 167 252
rect 118 203 122 207
rect 73 158 77 162
rect 28 113 32 117
rect 19 90 23 94
rect 34 96 38 100
rect 64 135 68 139
rect 79 141 83 145
rect 109 180 113 184
rect 124 186 128 190
rect 154 225 158 229
rect 169 231 173 235
rect 199 270 203 274
rect 214 276 218 280
rect 244 315 248 319
rect 259 321 263 325
rect 289 360 293 364
rect 304 366 308 370
rect 334 405 338 409
rect 349 411 353 415
rect 379 450 383 454
rect 394 456 398 460
rect 424 495 428 499
rect 439 501 443 505
rect 469 540 473 544
rect 484 546 488 550
rect 514 585 518 589
rect 529 591 533 595
rect 559 630 563 634
rect 574 636 578 640
rect 604 675 608 679
rect 619 681 623 685
rect 649 720 653 724
rect 664 726 668 730
rect 694 765 698 769
rect 709 771 713 775
rect 739 810 743 814
rect 754 816 758 820
rect 784 855 788 859
rect 799 861 803 865
rect 838 878 842 882
rect 793 833 797 837
rect 748 788 752 792
rect 703 743 707 747
rect 658 698 662 702
rect 613 653 617 657
rect 568 608 572 612
rect 523 563 527 567
rect 478 518 482 522
rect 433 473 437 477
rect 388 428 392 432
rect 343 383 347 387
rect 298 338 302 342
rect 253 293 257 297
rect 208 248 212 252
rect 163 203 167 207
rect 118 158 122 162
rect 73 113 77 117
rect 28 68 32 72
rect 19 45 23 49
rect 34 51 38 55
rect 64 90 68 94
rect 79 96 83 100
rect 109 135 113 139
rect 124 141 128 145
rect 154 180 158 184
rect 169 186 173 190
rect 199 225 203 229
rect 214 231 218 235
rect 244 270 248 274
rect 259 276 263 280
rect 289 315 293 319
rect 304 321 308 325
rect 334 360 338 364
rect 349 366 353 370
rect 379 405 383 409
rect 394 411 398 415
rect 424 450 428 454
rect 439 456 443 460
rect 469 495 473 499
rect 484 501 488 505
rect 514 540 518 544
rect 529 546 533 550
rect 559 585 563 589
rect 574 591 578 595
rect 604 630 608 634
rect 619 636 623 640
rect 649 675 653 679
rect 664 681 668 685
rect 694 720 698 724
rect 709 726 713 730
rect 739 765 743 769
rect 754 771 758 775
rect 784 810 788 814
rect 799 816 803 820
rect 829 855 833 859
rect 844 861 848 865
rect 883 878 887 882
rect 838 833 842 837
rect 793 788 797 792
rect 748 743 752 747
rect 703 698 707 702
rect 658 653 662 657
rect 613 608 617 612
rect 568 563 572 567
rect 523 518 527 522
rect 478 473 482 477
rect 433 428 437 432
rect 388 383 392 387
rect 343 338 347 342
rect 298 293 302 297
rect 253 248 257 252
rect 208 203 212 207
rect 163 158 167 162
rect 118 113 122 117
rect 73 68 77 72
rect 28 23 32 27
rect 19 0 23 4
rect 34 6 38 10
rect 64 45 68 49
rect 79 51 83 55
rect 109 90 113 94
rect 124 96 128 100
rect 154 135 158 139
rect 169 141 173 145
rect 199 180 203 184
rect 214 186 218 190
rect 244 225 248 229
rect 259 231 263 235
rect 289 270 293 274
rect 304 276 308 280
rect 334 315 338 319
rect 349 321 353 325
rect 379 360 383 364
rect 394 366 398 370
rect 424 405 428 409
rect 439 411 443 415
rect 469 450 473 454
rect 484 456 488 460
rect 514 495 518 499
rect 529 501 533 505
rect 559 540 563 544
rect 574 546 578 550
rect 604 585 608 589
rect 619 591 623 595
rect 649 630 653 634
rect 664 636 668 640
rect 694 675 698 679
rect 709 681 713 685
rect 739 720 743 724
rect 754 726 758 730
rect 784 765 788 769
rect 799 771 803 775
rect 829 810 833 814
rect 844 816 848 820
rect 874 855 878 859
rect 889 861 893 865
rect 883 833 887 837
rect 838 788 842 792
rect 793 743 797 747
rect 748 698 752 702
rect 703 653 707 657
rect 658 608 662 612
rect 613 563 617 567
rect 568 518 572 522
rect 523 473 527 477
rect 478 428 482 432
rect 433 383 437 387
rect 388 338 392 342
rect 343 293 347 297
rect 298 248 302 252
rect 253 203 257 207
rect 208 158 212 162
rect 163 113 167 117
rect 118 68 122 72
rect 73 23 77 27
rect 64 0 68 4
rect 79 6 83 10
rect 109 45 113 49
rect 124 51 128 55
rect 154 90 158 94
rect 169 96 173 100
rect 199 135 203 139
rect 214 141 218 145
rect 244 180 248 184
rect 259 186 263 190
rect 289 225 293 229
rect 304 231 308 235
rect 334 270 338 274
rect 349 276 353 280
rect 379 315 383 319
rect 394 321 398 325
rect 424 360 428 364
rect 439 366 443 370
rect 469 405 473 409
rect 484 411 488 415
rect 514 450 518 454
rect 529 456 533 460
rect 559 495 563 499
rect 574 501 578 505
rect 604 540 608 544
rect 619 546 623 550
rect 649 585 653 589
rect 664 591 668 595
rect 694 630 698 634
rect 709 636 713 640
rect 739 675 743 679
rect 754 681 758 685
rect 784 720 788 724
rect 799 726 803 730
rect 829 765 833 769
rect 844 771 848 775
rect 874 810 878 814
rect 889 816 893 820
rect 883 788 887 792
rect 838 743 842 747
rect 793 698 797 702
rect 748 653 752 657
rect 703 608 707 612
rect 658 563 662 567
rect 613 518 617 522
rect 568 473 572 477
rect 523 428 527 432
rect 478 383 482 387
rect 433 338 437 342
rect 388 293 392 297
rect 343 248 347 252
rect 298 203 302 207
rect 253 158 257 162
rect 208 113 212 117
rect 163 68 167 72
rect 118 23 122 27
rect 109 0 113 4
rect 124 6 128 10
rect 154 45 158 49
rect 169 51 173 55
rect 199 90 203 94
rect 214 96 218 100
rect 244 135 248 139
rect 259 141 263 145
rect 289 180 293 184
rect 304 186 308 190
rect 334 225 338 229
rect 349 231 353 235
rect 379 270 383 274
rect 394 276 398 280
rect 424 315 428 319
rect 439 321 443 325
rect 469 360 473 364
rect 484 366 488 370
rect 514 405 518 409
rect 529 411 533 415
rect 559 450 563 454
rect 574 456 578 460
rect 604 495 608 499
rect 619 501 623 505
rect 649 540 653 544
rect 664 546 668 550
rect 694 585 698 589
rect 709 591 713 595
rect 739 630 743 634
rect 754 636 758 640
rect 784 675 788 679
rect 799 681 803 685
rect 829 720 833 724
rect 844 726 848 730
rect 874 765 878 769
rect 889 771 893 775
rect 883 743 887 747
rect 838 698 842 702
rect 793 653 797 657
rect 748 608 752 612
rect 703 563 707 567
rect 658 518 662 522
rect 613 473 617 477
rect 568 428 572 432
rect 523 383 527 387
rect 478 338 482 342
rect 433 293 437 297
rect 388 248 392 252
rect 343 203 347 207
rect 298 158 302 162
rect 253 113 257 117
rect 208 68 212 72
rect 163 23 167 27
rect 154 0 158 4
rect 169 6 173 10
rect 199 45 203 49
rect 214 51 218 55
rect 244 90 248 94
rect 259 96 263 100
rect 289 135 293 139
rect 304 141 308 145
rect 334 180 338 184
rect 349 186 353 190
rect 379 225 383 229
rect 394 231 398 235
rect 424 270 428 274
rect 439 276 443 280
rect 469 315 473 319
rect 484 321 488 325
rect 514 360 518 364
rect 529 366 533 370
rect 559 405 563 409
rect 574 411 578 415
rect 604 450 608 454
rect 619 456 623 460
rect 649 495 653 499
rect 664 501 668 505
rect 694 540 698 544
rect 709 546 713 550
rect 739 585 743 589
rect 754 591 758 595
rect 784 630 788 634
rect 799 636 803 640
rect 829 675 833 679
rect 844 681 848 685
rect 874 720 878 724
rect 889 726 893 730
rect 883 698 887 702
rect 838 653 842 657
rect 793 608 797 612
rect 748 563 752 567
rect 703 518 707 522
rect 658 473 662 477
rect 613 428 617 432
rect 568 383 572 387
rect 523 338 527 342
rect 478 293 482 297
rect 433 248 437 252
rect 388 203 392 207
rect 343 158 347 162
rect 298 113 302 117
rect 253 68 257 72
rect 208 23 212 27
rect 199 0 203 4
rect 214 6 218 10
rect 244 45 248 49
rect 259 51 263 55
rect 289 90 293 94
rect 304 96 308 100
rect 334 135 338 139
rect 349 141 353 145
rect 379 180 383 184
rect 394 186 398 190
rect 424 225 428 229
rect 439 231 443 235
rect 469 270 473 274
rect 484 276 488 280
rect 514 315 518 319
rect 529 321 533 325
rect 559 360 563 364
rect 574 366 578 370
rect 604 405 608 409
rect 619 411 623 415
rect 649 450 653 454
rect 664 456 668 460
rect 694 495 698 499
rect 709 501 713 505
rect 739 540 743 544
rect 754 546 758 550
rect 784 585 788 589
rect 799 591 803 595
rect 829 630 833 634
rect 844 636 848 640
rect 874 675 878 679
rect 889 681 893 685
rect 883 653 887 657
rect 838 608 842 612
rect 793 563 797 567
rect 748 518 752 522
rect 703 473 707 477
rect 658 428 662 432
rect 613 383 617 387
rect 568 338 572 342
rect 523 293 527 297
rect 478 248 482 252
rect 433 203 437 207
rect 388 158 392 162
rect 343 113 347 117
rect 298 68 302 72
rect 253 23 257 27
rect 244 0 248 4
rect 259 6 263 10
rect 289 45 293 49
rect 304 51 308 55
rect 334 90 338 94
rect 349 96 353 100
rect 379 135 383 139
rect 394 141 398 145
rect 424 180 428 184
rect 439 186 443 190
rect 469 225 473 229
rect 484 231 488 235
rect 514 270 518 274
rect 529 276 533 280
rect 559 315 563 319
rect 574 321 578 325
rect 604 360 608 364
rect 619 366 623 370
rect 649 405 653 409
rect 664 411 668 415
rect 694 450 698 454
rect 709 456 713 460
rect 739 495 743 499
rect 754 501 758 505
rect 784 540 788 544
rect 799 546 803 550
rect 829 585 833 589
rect 844 591 848 595
rect 874 630 878 634
rect 889 636 893 640
rect 883 608 887 612
rect 838 563 842 567
rect 793 518 797 522
rect 748 473 752 477
rect 703 428 707 432
rect 658 383 662 387
rect 613 338 617 342
rect 568 293 572 297
rect 523 248 527 252
rect 478 203 482 207
rect 433 158 437 162
rect 388 113 392 117
rect 343 68 347 72
rect 298 23 302 27
rect 289 0 293 4
rect 304 6 308 10
rect 334 45 338 49
rect 349 51 353 55
rect 379 90 383 94
rect 394 96 398 100
rect 424 135 428 139
rect 439 141 443 145
rect 469 180 473 184
rect 484 186 488 190
rect 514 225 518 229
rect 529 231 533 235
rect 559 270 563 274
rect 574 276 578 280
rect 604 315 608 319
rect 619 321 623 325
rect 649 360 653 364
rect 664 366 668 370
rect 694 405 698 409
rect 709 411 713 415
rect 739 450 743 454
rect 754 456 758 460
rect 784 495 788 499
rect 799 501 803 505
rect 829 540 833 544
rect 844 546 848 550
rect 874 585 878 589
rect 889 591 893 595
rect 883 563 887 567
rect 838 518 842 522
rect 793 473 797 477
rect 748 428 752 432
rect 703 383 707 387
rect 658 338 662 342
rect 613 293 617 297
rect 568 248 572 252
rect 523 203 527 207
rect 478 158 482 162
rect 433 113 437 117
rect 388 68 392 72
rect 343 23 347 27
rect 334 0 338 4
rect 349 6 353 10
rect 379 45 383 49
rect 394 51 398 55
rect 424 90 428 94
rect 439 96 443 100
rect 469 135 473 139
rect 484 141 488 145
rect 514 180 518 184
rect 529 186 533 190
rect 559 225 563 229
rect 574 231 578 235
rect 604 270 608 274
rect 619 276 623 280
rect 649 315 653 319
rect 664 321 668 325
rect 694 360 698 364
rect 709 366 713 370
rect 739 405 743 409
rect 754 411 758 415
rect 784 450 788 454
rect 799 456 803 460
rect 829 495 833 499
rect 844 501 848 505
rect 874 540 878 544
rect 889 546 893 550
rect 883 518 887 522
rect 838 473 842 477
rect 793 428 797 432
rect 748 383 752 387
rect 703 338 707 342
rect 658 293 662 297
rect 613 248 617 252
rect 568 203 572 207
rect 523 158 527 162
rect 478 113 482 117
rect 433 68 437 72
rect 388 23 392 27
rect 379 0 383 4
rect 394 6 398 10
rect 424 45 428 49
rect 439 51 443 55
rect 469 90 473 94
rect 484 96 488 100
rect 514 135 518 139
rect 529 141 533 145
rect 559 180 563 184
rect 574 186 578 190
rect 604 225 608 229
rect 619 231 623 235
rect 649 270 653 274
rect 664 276 668 280
rect 694 315 698 319
rect 709 321 713 325
rect 739 360 743 364
rect 754 366 758 370
rect 784 405 788 409
rect 799 411 803 415
rect 829 450 833 454
rect 844 456 848 460
rect 874 495 878 499
rect 889 501 893 505
rect 883 473 887 477
rect 838 428 842 432
rect 793 383 797 387
rect 748 338 752 342
rect 703 293 707 297
rect 658 248 662 252
rect 613 203 617 207
rect 568 158 572 162
rect 523 113 527 117
rect 478 68 482 72
rect 433 23 437 27
rect 424 0 428 4
rect 439 6 443 10
rect 469 45 473 49
rect 484 51 488 55
rect 514 90 518 94
rect 529 96 533 100
rect 559 135 563 139
rect 574 141 578 145
rect 604 180 608 184
rect 619 186 623 190
rect 649 225 653 229
rect 664 231 668 235
rect 694 270 698 274
rect 709 276 713 280
rect 739 315 743 319
rect 754 321 758 325
rect 784 360 788 364
rect 799 366 803 370
rect 829 405 833 409
rect 844 411 848 415
rect 874 450 878 454
rect 889 456 893 460
rect 883 428 887 432
rect 838 383 842 387
rect 793 338 797 342
rect 748 293 752 297
rect 703 248 707 252
rect 658 203 662 207
rect 613 158 617 162
rect 568 113 572 117
rect 523 68 527 72
rect 478 23 482 27
rect 469 0 473 4
rect 484 6 488 10
rect 514 45 518 49
rect 529 51 533 55
rect 559 90 563 94
rect 574 96 578 100
rect 604 135 608 139
rect 619 141 623 145
rect 649 180 653 184
rect 664 186 668 190
rect 694 225 698 229
rect 709 231 713 235
rect 739 270 743 274
rect 754 276 758 280
rect 784 315 788 319
rect 799 321 803 325
rect 829 360 833 364
rect 844 366 848 370
rect 874 405 878 409
rect 889 411 893 415
rect 883 383 887 387
rect 838 338 842 342
rect 793 293 797 297
rect 748 248 752 252
rect 703 203 707 207
rect 658 158 662 162
rect 613 113 617 117
rect 568 68 572 72
rect 523 23 527 27
rect 514 0 518 4
rect 529 6 533 10
rect 559 45 563 49
rect 574 51 578 55
rect 604 90 608 94
rect 619 96 623 100
rect 649 135 653 139
rect 664 141 668 145
rect 694 180 698 184
rect 709 186 713 190
rect 739 225 743 229
rect 754 231 758 235
rect 784 270 788 274
rect 799 276 803 280
rect 829 315 833 319
rect 844 321 848 325
rect 874 360 878 364
rect 889 366 893 370
rect 883 338 887 342
rect 838 293 842 297
rect 793 248 797 252
rect 748 203 752 207
rect 703 158 707 162
rect 658 113 662 117
rect 613 68 617 72
rect 568 23 572 27
rect 559 0 563 4
rect 574 6 578 10
rect 604 45 608 49
rect 619 51 623 55
rect 649 90 653 94
rect 664 96 668 100
rect 694 135 698 139
rect 709 141 713 145
rect 739 180 743 184
rect 754 186 758 190
rect 784 225 788 229
rect 799 231 803 235
rect 829 270 833 274
rect 844 276 848 280
rect 874 315 878 319
rect 889 321 893 325
rect 883 293 887 297
rect 838 248 842 252
rect 793 203 797 207
rect 748 158 752 162
rect 703 113 707 117
rect 658 68 662 72
rect 613 23 617 27
rect 604 0 608 4
rect 619 6 623 10
rect 649 45 653 49
rect 664 51 668 55
rect 694 90 698 94
rect 709 96 713 100
rect 739 135 743 139
rect 754 141 758 145
rect 784 180 788 184
rect 799 186 803 190
rect 829 225 833 229
rect 844 231 848 235
rect 874 270 878 274
rect 889 276 893 280
rect 883 248 887 252
rect 838 203 842 207
rect 793 158 797 162
rect 748 113 752 117
rect 703 68 707 72
rect 658 23 662 27
rect 649 0 653 4
rect 664 6 668 10
rect 694 45 698 49
rect 709 51 713 55
rect 739 90 743 94
rect 754 96 758 100
rect 784 135 788 139
rect 799 141 803 145
rect 829 180 833 184
rect 844 186 848 190
rect 874 225 878 229
rect 889 231 893 235
rect 883 203 887 207
rect 838 158 842 162
rect 793 113 797 117
rect 748 68 752 72
rect 703 23 707 27
rect 694 0 698 4
rect 709 6 713 10
rect 739 45 743 49
rect 754 51 758 55
rect 784 90 788 94
rect 799 96 803 100
rect 829 135 833 139
rect 844 141 848 145
rect 874 180 878 184
rect 889 186 893 190
rect 883 158 887 162
rect 838 113 842 117
rect 793 68 797 72
rect 748 23 752 27
rect 739 0 743 4
rect 754 6 758 10
rect 784 45 788 49
rect 799 51 803 55
rect 829 90 833 94
rect 844 96 848 100
rect 874 135 878 139
rect 889 141 893 145
rect 883 113 887 117
rect 838 68 842 72
rect 793 23 797 27
rect 784 0 788 4
rect 799 6 803 10
rect 829 45 833 49
rect 844 51 848 55
rect 874 90 878 94
rect 889 96 893 100
rect 883 68 887 72
rect 838 23 842 27
rect 829 0 833 4
rect 844 6 848 10
rect 874 45 878 49
rect 889 51 893 55
rect 883 23 887 27
rect 874 0 878 4
rect 889 6 893 10
rect -300 -161 -296 -157
rect -277 -169 -273 -165
rect -282 -176 -278 -172
rect -188 -158 -184 -154
rect -257 -179 -253 -175
rect -197 -181 -193 -177
rect -182 -175 -178 -171
<< metal2 >>
rect 0 879 28 882
rect 32 879 73 882
rect 77 879 118 882
rect 122 879 163 882
rect 167 879 208 882
rect 212 879 253 882
rect 257 879 298 882
rect 302 879 343 882
rect 347 879 388 882
rect 392 879 433 882
rect 437 879 478 882
rect 482 879 523 882
rect 527 879 568 882
rect 572 879 613 882
rect 617 879 658 882
rect 662 879 703 882
rect 707 879 748 882
rect 752 879 793 882
rect 797 879 838 882
rect 842 879 883 882
rect 887 879 900 882
rect 0 862 34 865
rect 38 862 79 865
rect 83 862 124 865
rect 128 862 169 865
rect 173 862 214 865
rect 218 862 259 865
rect 263 862 304 865
rect 308 862 349 865
rect 353 862 394 865
rect 398 862 439 865
rect 443 862 484 865
rect 488 862 529 865
rect 533 862 574 865
rect 578 862 619 865
rect 623 862 664 865
rect 668 862 709 865
rect 713 862 754 865
rect 758 862 799 865
rect 803 862 844 865
rect 848 862 889 865
rect 893 862 900 865
rect 0 855 19 858
rect 23 855 64 858
rect 68 855 109 858
rect 113 855 154 858
rect 158 855 199 858
rect 203 855 244 858
rect 248 855 289 858
rect 293 855 334 858
rect 338 855 379 858
rect 383 855 424 858
rect 428 855 469 858
rect 473 855 514 858
rect 518 855 559 858
rect 563 855 604 858
rect 608 855 649 858
rect 653 855 694 858
rect 698 855 739 858
rect 743 855 784 858
rect 788 855 829 858
rect 833 855 874 858
rect 878 855 900 858
rect 0 834 28 837
rect 32 834 73 837
rect 77 834 118 837
rect 122 834 163 837
rect 167 834 208 837
rect 212 834 253 837
rect 257 834 298 837
rect 302 834 343 837
rect 347 834 388 837
rect 392 834 433 837
rect 437 834 478 837
rect 482 834 523 837
rect 527 834 568 837
rect 572 834 613 837
rect 617 834 658 837
rect 662 834 703 837
rect 707 834 748 837
rect 752 834 793 837
rect 797 834 838 837
rect 842 834 883 837
rect 887 834 900 837
rect 0 817 34 820
rect 38 817 79 820
rect 83 817 124 820
rect 128 817 169 820
rect 173 817 214 820
rect 218 817 259 820
rect 263 817 304 820
rect 308 817 349 820
rect 353 817 394 820
rect 398 817 439 820
rect 443 817 484 820
rect 488 817 529 820
rect 533 817 574 820
rect 578 817 619 820
rect 623 817 664 820
rect 668 817 709 820
rect 713 817 754 820
rect 758 817 799 820
rect 803 817 844 820
rect 848 817 889 820
rect 893 817 900 820
rect 0 810 19 813
rect 23 810 64 813
rect 68 810 109 813
rect 113 810 154 813
rect 158 810 199 813
rect 203 810 244 813
rect 248 810 289 813
rect 293 810 334 813
rect 338 810 379 813
rect 383 810 424 813
rect 428 810 469 813
rect 473 810 514 813
rect 518 810 559 813
rect 563 810 604 813
rect 608 810 649 813
rect 653 810 694 813
rect 698 810 739 813
rect 743 810 784 813
rect 788 810 829 813
rect 833 810 874 813
rect 878 810 900 813
rect 0 789 28 792
rect 32 789 73 792
rect 77 789 118 792
rect 122 789 163 792
rect 167 789 208 792
rect 212 789 253 792
rect 257 789 298 792
rect 302 789 343 792
rect 347 789 388 792
rect 392 789 433 792
rect 437 789 478 792
rect 482 789 523 792
rect 527 789 568 792
rect 572 789 613 792
rect 617 789 658 792
rect 662 789 703 792
rect 707 789 748 792
rect 752 789 793 792
rect 797 789 838 792
rect 842 789 883 792
rect 887 789 900 792
rect 0 772 34 775
rect 38 772 79 775
rect 83 772 124 775
rect 128 772 169 775
rect 173 772 214 775
rect 218 772 259 775
rect 263 772 304 775
rect 308 772 349 775
rect 353 772 394 775
rect 398 772 439 775
rect 443 772 484 775
rect 488 772 529 775
rect 533 772 574 775
rect 578 772 619 775
rect 623 772 664 775
rect 668 772 709 775
rect 713 772 754 775
rect 758 772 799 775
rect 803 772 844 775
rect 848 772 889 775
rect 893 772 900 775
rect 0 765 19 768
rect 23 765 64 768
rect 68 765 109 768
rect 113 765 154 768
rect 158 765 199 768
rect 203 765 244 768
rect 248 765 289 768
rect 293 765 334 768
rect 338 765 379 768
rect 383 765 424 768
rect 428 765 469 768
rect 473 765 514 768
rect 518 765 559 768
rect 563 765 604 768
rect 608 765 649 768
rect 653 765 694 768
rect 698 765 739 768
rect 743 765 784 768
rect 788 765 829 768
rect 833 765 874 768
rect 878 765 900 768
rect 0 744 28 747
rect 32 744 73 747
rect 77 744 118 747
rect 122 744 163 747
rect 167 744 208 747
rect 212 744 253 747
rect 257 744 298 747
rect 302 744 343 747
rect 347 744 388 747
rect 392 744 433 747
rect 437 744 478 747
rect 482 744 523 747
rect 527 744 568 747
rect 572 744 613 747
rect 617 744 658 747
rect 662 744 703 747
rect 707 744 748 747
rect 752 744 793 747
rect 797 744 838 747
rect 842 744 883 747
rect 887 744 900 747
rect 0 727 34 730
rect 38 727 79 730
rect 83 727 124 730
rect 128 727 169 730
rect 173 727 214 730
rect 218 727 259 730
rect 263 727 304 730
rect 308 727 349 730
rect 353 727 394 730
rect 398 727 439 730
rect 443 727 484 730
rect 488 727 529 730
rect 533 727 574 730
rect 578 727 619 730
rect 623 727 664 730
rect 668 727 709 730
rect 713 727 754 730
rect 758 727 799 730
rect 803 727 844 730
rect 848 727 889 730
rect 893 727 900 730
rect 0 720 19 723
rect 23 720 64 723
rect 68 720 109 723
rect 113 720 154 723
rect 158 720 199 723
rect 203 720 244 723
rect 248 720 289 723
rect 293 720 334 723
rect 338 720 379 723
rect 383 720 424 723
rect 428 720 469 723
rect 473 720 514 723
rect 518 720 559 723
rect 563 720 604 723
rect 608 720 649 723
rect 653 720 694 723
rect 698 720 739 723
rect 743 720 784 723
rect 788 720 829 723
rect 833 720 874 723
rect 878 720 900 723
rect 0 699 28 702
rect 32 699 73 702
rect 77 699 118 702
rect 122 699 163 702
rect 167 699 208 702
rect 212 699 253 702
rect 257 699 298 702
rect 302 699 343 702
rect 347 699 388 702
rect 392 699 433 702
rect 437 699 478 702
rect 482 699 523 702
rect 527 699 568 702
rect 572 699 613 702
rect 617 699 658 702
rect 662 699 703 702
rect 707 699 748 702
rect 752 699 793 702
rect 797 699 838 702
rect 842 699 883 702
rect 887 699 900 702
rect 0 682 34 685
rect 38 682 79 685
rect 83 682 124 685
rect 128 682 169 685
rect 173 682 214 685
rect 218 682 259 685
rect 263 682 304 685
rect 308 682 349 685
rect 353 682 394 685
rect 398 682 439 685
rect 443 682 484 685
rect 488 682 529 685
rect 533 682 574 685
rect 578 682 619 685
rect 623 682 664 685
rect 668 682 709 685
rect 713 682 754 685
rect 758 682 799 685
rect 803 682 844 685
rect 848 682 889 685
rect 893 682 900 685
rect 0 675 19 678
rect 23 675 64 678
rect 68 675 109 678
rect 113 675 154 678
rect 158 675 199 678
rect 203 675 244 678
rect 248 675 289 678
rect 293 675 334 678
rect 338 675 379 678
rect 383 675 424 678
rect 428 675 469 678
rect 473 675 514 678
rect 518 675 559 678
rect 563 675 604 678
rect 608 675 649 678
rect 653 675 694 678
rect 698 675 739 678
rect 743 675 784 678
rect 788 675 829 678
rect 833 675 874 678
rect 878 675 900 678
rect 0 654 28 657
rect 32 654 73 657
rect 77 654 118 657
rect 122 654 163 657
rect 167 654 208 657
rect 212 654 253 657
rect 257 654 298 657
rect 302 654 343 657
rect 347 654 388 657
rect 392 654 433 657
rect 437 654 478 657
rect 482 654 523 657
rect 527 654 568 657
rect 572 654 613 657
rect 617 654 658 657
rect 662 654 703 657
rect 707 654 748 657
rect 752 654 793 657
rect 797 654 838 657
rect 842 654 883 657
rect 887 654 900 657
rect 0 637 34 640
rect 38 637 79 640
rect 83 637 124 640
rect 128 637 169 640
rect 173 637 214 640
rect 218 637 259 640
rect 263 637 304 640
rect 308 637 349 640
rect 353 637 394 640
rect 398 637 439 640
rect 443 637 484 640
rect 488 637 529 640
rect 533 637 574 640
rect 578 637 619 640
rect 623 637 664 640
rect 668 637 709 640
rect 713 637 754 640
rect 758 637 799 640
rect 803 637 844 640
rect 848 637 889 640
rect 893 637 900 640
rect 0 630 19 633
rect 23 630 64 633
rect 68 630 109 633
rect 113 630 154 633
rect 158 630 199 633
rect 203 630 244 633
rect 248 630 289 633
rect 293 630 334 633
rect 338 630 379 633
rect 383 630 424 633
rect 428 630 469 633
rect 473 630 514 633
rect 518 630 559 633
rect 563 630 604 633
rect 608 630 649 633
rect 653 630 694 633
rect 698 630 739 633
rect 743 630 784 633
rect 788 630 829 633
rect 833 630 874 633
rect 878 630 900 633
rect 0 609 28 612
rect 32 609 73 612
rect 77 609 118 612
rect 122 609 163 612
rect 167 609 208 612
rect 212 609 253 612
rect 257 609 298 612
rect 302 609 343 612
rect 347 609 388 612
rect 392 609 433 612
rect 437 609 478 612
rect 482 609 523 612
rect 527 609 568 612
rect 572 609 613 612
rect 617 609 658 612
rect 662 609 703 612
rect 707 609 748 612
rect 752 609 793 612
rect 797 609 838 612
rect 842 609 883 612
rect 887 609 900 612
rect 0 592 34 595
rect 38 592 79 595
rect 83 592 124 595
rect 128 592 169 595
rect 173 592 214 595
rect 218 592 259 595
rect 263 592 304 595
rect 308 592 349 595
rect 353 592 394 595
rect 398 592 439 595
rect 443 592 484 595
rect 488 592 529 595
rect 533 592 574 595
rect 578 592 619 595
rect 623 592 664 595
rect 668 592 709 595
rect 713 592 754 595
rect 758 592 799 595
rect 803 592 844 595
rect 848 592 889 595
rect 893 592 900 595
rect 0 585 19 588
rect 23 585 64 588
rect 68 585 109 588
rect 113 585 154 588
rect 158 585 199 588
rect 203 585 244 588
rect 248 585 289 588
rect 293 585 334 588
rect 338 585 379 588
rect 383 585 424 588
rect 428 585 469 588
rect 473 585 514 588
rect 518 585 559 588
rect 563 585 604 588
rect 608 585 649 588
rect 653 585 694 588
rect 698 585 739 588
rect 743 585 784 588
rect 788 585 829 588
rect 833 585 874 588
rect 878 585 900 588
rect 0 564 28 567
rect 32 564 73 567
rect 77 564 118 567
rect 122 564 163 567
rect 167 564 208 567
rect 212 564 253 567
rect 257 564 298 567
rect 302 564 343 567
rect 347 564 388 567
rect 392 564 433 567
rect 437 564 478 567
rect 482 564 523 567
rect 527 564 568 567
rect 572 564 613 567
rect 617 564 658 567
rect 662 564 703 567
rect 707 564 748 567
rect 752 564 793 567
rect 797 564 838 567
rect 842 564 883 567
rect 887 564 900 567
rect 0 547 34 550
rect 38 547 79 550
rect 83 547 124 550
rect 128 547 169 550
rect 173 547 214 550
rect 218 547 259 550
rect 263 547 304 550
rect 308 547 349 550
rect 353 547 394 550
rect 398 547 439 550
rect 443 547 484 550
rect 488 547 529 550
rect 533 547 574 550
rect 578 547 619 550
rect 623 547 664 550
rect 668 547 709 550
rect 713 547 754 550
rect 758 547 799 550
rect 803 547 844 550
rect 848 547 889 550
rect 893 547 900 550
rect 0 540 19 543
rect 23 540 64 543
rect 68 540 109 543
rect 113 540 154 543
rect 158 540 199 543
rect 203 540 244 543
rect 248 540 289 543
rect 293 540 334 543
rect 338 540 379 543
rect 383 540 424 543
rect 428 540 469 543
rect 473 540 514 543
rect 518 540 559 543
rect 563 540 604 543
rect 608 540 649 543
rect 653 540 694 543
rect 698 540 739 543
rect 743 540 784 543
rect 788 540 829 543
rect 833 540 874 543
rect 878 540 900 543
rect 0 519 28 522
rect 32 519 73 522
rect 77 519 118 522
rect 122 519 163 522
rect 167 519 208 522
rect 212 519 253 522
rect 257 519 298 522
rect 302 519 343 522
rect 347 519 388 522
rect 392 519 433 522
rect 437 519 478 522
rect 482 519 523 522
rect 527 519 568 522
rect 572 519 613 522
rect 617 519 658 522
rect 662 519 703 522
rect 707 519 748 522
rect 752 519 793 522
rect 797 519 838 522
rect 842 519 883 522
rect 887 519 900 522
rect 0 502 34 505
rect 38 502 79 505
rect 83 502 124 505
rect 128 502 169 505
rect 173 502 214 505
rect 218 502 259 505
rect 263 502 304 505
rect 308 502 349 505
rect 353 502 394 505
rect 398 502 439 505
rect 443 502 484 505
rect 488 502 529 505
rect 533 502 574 505
rect 578 502 619 505
rect 623 502 664 505
rect 668 502 709 505
rect 713 502 754 505
rect 758 502 799 505
rect 803 502 844 505
rect 848 502 889 505
rect 893 502 900 505
rect 0 495 19 498
rect 23 495 64 498
rect 68 495 109 498
rect 113 495 154 498
rect 158 495 199 498
rect 203 495 244 498
rect 248 495 289 498
rect 293 495 334 498
rect 338 495 379 498
rect 383 495 424 498
rect 428 495 469 498
rect 473 495 514 498
rect 518 495 559 498
rect 563 495 604 498
rect 608 495 649 498
rect 653 495 694 498
rect 698 495 739 498
rect 743 495 784 498
rect 788 495 829 498
rect 833 495 874 498
rect 878 495 900 498
rect 0 474 28 477
rect 32 474 73 477
rect 77 474 118 477
rect 122 474 163 477
rect 167 474 208 477
rect 212 474 253 477
rect 257 474 298 477
rect 302 474 343 477
rect 347 474 388 477
rect 392 474 433 477
rect 437 474 478 477
rect 482 474 523 477
rect 527 474 568 477
rect 572 474 613 477
rect 617 474 658 477
rect 662 474 703 477
rect 707 474 748 477
rect 752 474 793 477
rect 797 474 838 477
rect 842 474 883 477
rect 887 474 900 477
rect 0 457 34 460
rect 38 457 79 460
rect 83 457 124 460
rect 128 457 169 460
rect 173 457 214 460
rect 218 457 259 460
rect 263 457 304 460
rect 308 457 349 460
rect 353 457 394 460
rect 398 457 439 460
rect 443 457 484 460
rect 488 457 529 460
rect 533 457 574 460
rect 578 457 619 460
rect 623 457 664 460
rect 668 457 709 460
rect 713 457 754 460
rect 758 457 799 460
rect 803 457 844 460
rect 848 457 889 460
rect 893 457 900 460
rect 0 450 19 453
rect 23 450 64 453
rect 68 450 109 453
rect 113 450 154 453
rect 158 450 199 453
rect 203 450 244 453
rect 248 450 289 453
rect 293 450 334 453
rect 338 450 379 453
rect 383 450 424 453
rect 428 450 469 453
rect 473 450 514 453
rect 518 450 559 453
rect 563 450 604 453
rect 608 450 649 453
rect 653 450 694 453
rect 698 450 739 453
rect 743 450 784 453
rect 788 450 829 453
rect 833 450 874 453
rect 878 450 900 453
rect 0 429 28 432
rect 32 429 73 432
rect 77 429 118 432
rect 122 429 163 432
rect 167 429 208 432
rect 212 429 253 432
rect 257 429 298 432
rect 302 429 343 432
rect 347 429 388 432
rect 392 429 433 432
rect 437 429 478 432
rect 482 429 523 432
rect 527 429 568 432
rect 572 429 613 432
rect 617 429 658 432
rect 662 429 703 432
rect 707 429 748 432
rect 752 429 793 432
rect 797 429 838 432
rect 842 429 883 432
rect 887 429 900 432
rect 0 412 34 415
rect 38 412 79 415
rect 83 412 124 415
rect 128 412 169 415
rect 173 412 214 415
rect 218 412 259 415
rect 263 412 304 415
rect 308 412 349 415
rect 353 412 394 415
rect 398 412 439 415
rect 443 412 484 415
rect 488 412 529 415
rect 533 412 574 415
rect 578 412 619 415
rect 623 412 664 415
rect 668 412 709 415
rect 713 412 754 415
rect 758 412 799 415
rect 803 412 844 415
rect 848 412 889 415
rect 893 412 900 415
rect 0 405 19 408
rect 23 405 64 408
rect 68 405 109 408
rect 113 405 154 408
rect 158 405 199 408
rect 203 405 244 408
rect 248 405 289 408
rect 293 405 334 408
rect 338 405 379 408
rect 383 405 424 408
rect 428 405 469 408
rect 473 405 514 408
rect 518 405 559 408
rect 563 405 604 408
rect 608 405 649 408
rect 653 405 694 408
rect 698 405 739 408
rect 743 405 784 408
rect 788 405 829 408
rect 833 405 874 408
rect 878 405 900 408
rect 0 384 28 387
rect 32 384 73 387
rect 77 384 118 387
rect 122 384 163 387
rect 167 384 208 387
rect 212 384 253 387
rect 257 384 298 387
rect 302 384 343 387
rect 347 384 388 387
rect 392 384 433 387
rect 437 384 478 387
rect 482 384 523 387
rect 527 384 568 387
rect 572 384 613 387
rect 617 384 658 387
rect 662 384 703 387
rect 707 384 748 387
rect 752 384 793 387
rect 797 384 838 387
rect 842 384 883 387
rect 887 384 900 387
rect 0 367 34 370
rect 38 367 79 370
rect 83 367 124 370
rect 128 367 169 370
rect 173 367 214 370
rect 218 367 259 370
rect 263 367 304 370
rect 308 367 349 370
rect 353 367 394 370
rect 398 367 439 370
rect 443 367 484 370
rect 488 367 529 370
rect 533 367 574 370
rect 578 367 619 370
rect 623 367 664 370
rect 668 367 709 370
rect 713 367 754 370
rect 758 367 799 370
rect 803 367 844 370
rect 848 367 889 370
rect 893 367 900 370
rect 0 360 19 363
rect 23 360 64 363
rect 68 360 109 363
rect 113 360 154 363
rect 158 360 199 363
rect 203 360 244 363
rect 248 360 289 363
rect 293 360 334 363
rect 338 360 379 363
rect 383 360 424 363
rect 428 360 469 363
rect 473 360 514 363
rect 518 360 559 363
rect 563 360 604 363
rect 608 360 649 363
rect 653 360 694 363
rect 698 360 739 363
rect 743 360 784 363
rect 788 360 829 363
rect 833 360 874 363
rect 878 360 900 363
rect 0 339 28 342
rect 32 339 73 342
rect 77 339 118 342
rect 122 339 163 342
rect 167 339 208 342
rect 212 339 253 342
rect 257 339 298 342
rect 302 339 343 342
rect 347 339 388 342
rect 392 339 433 342
rect 437 339 478 342
rect 482 339 523 342
rect 527 339 568 342
rect 572 339 613 342
rect 617 339 658 342
rect 662 339 703 342
rect 707 339 748 342
rect 752 339 793 342
rect 797 339 838 342
rect 842 339 883 342
rect 887 339 900 342
rect 0 322 34 325
rect 38 322 79 325
rect 83 322 124 325
rect 128 322 169 325
rect 173 322 214 325
rect 218 322 259 325
rect 263 322 304 325
rect 308 322 349 325
rect 353 322 394 325
rect 398 322 439 325
rect 443 322 484 325
rect 488 322 529 325
rect 533 322 574 325
rect 578 322 619 325
rect 623 322 664 325
rect 668 322 709 325
rect 713 322 754 325
rect 758 322 799 325
rect 803 322 844 325
rect 848 322 889 325
rect 893 322 900 325
rect 0 315 19 318
rect 23 315 64 318
rect 68 315 109 318
rect 113 315 154 318
rect 158 315 199 318
rect 203 315 244 318
rect 248 315 289 318
rect 293 315 334 318
rect 338 315 379 318
rect 383 315 424 318
rect 428 315 469 318
rect 473 315 514 318
rect 518 315 559 318
rect 563 315 604 318
rect 608 315 649 318
rect 653 315 694 318
rect 698 315 739 318
rect 743 315 784 318
rect 788 315 829 318
rect 833 315 874 318
rect 878 315 900 318
rect 0 294 28 297
rect 32 294 73 297
rect 77 294 118 297
rect 122 294 163 297
rect 167 294 208 297
rect 212 294 253 297
rect 257 294 298 297
rect 302 294 343 297
rect 347 294 388 297
rect 392 294 433 297
rect 437 294 478 297
rect 482 294 523 297
rect 527 294 568 297
rect 572 294 613 297
rect 617 294 658 297
rect 662 294 703 297
rect 707 294 748 297
rect 752 294 793 297
rect 797 294 838 297
rect 842 294 883 297
rect 887 294 900 297
rect 0 277 34 280
rect 38 277 79 280
rect 83 277 124 280
rect 128 277 169 280
rect 173 277 214 280
rect 218 277 259 280
rect 263 277 304 280
rect 308 277 349 280
rect 353 277 394 280
rect 398 277 439 280
rect 443 277 484 280
rect 488 277 529 280
rect 533 277 574 280
rect 578 277 619 280
rect 623 277 664 280
rect 668 277 709 280
rect 713 277 754 280
rect 758 277 799 280
rect 803 277 844 280
rect 848 277 889 280
rect 893 277 900 280
rect 0 270 19 273
rect 23 270 64 273
rect 68 270 109 273
rect 113 270 154 273
rect 158 270 199 273
rect 203 270 244 273
rect 248 270 289 273
rect 293 270 334 273
rect 338 270 379 273
rect 383 270 424 273
rect 428 270 469 273
rect 473 270 514 273
rect 518 270 559 273
rect 563 270 604 273
rect 608 270 649 273
rect 653 270 694 273
rect 698 270 739 273
rect 743 270 784 273
rect 788 270 829 273
rect 833 270 874 273
rect 878 270 900 273
rect 0 249 28 252
rect 32 249 73 252
rect 77 249 118 252
rect 122 249 163 252
rect 167 249 208 252
rect 212 249 253 252
rect 257 249 298 252
rect 302 249 343 252
rect 347 249 388 252
rect 392 249 433 252
rect 437 249 478 252
rect 482 249 523 252
rect 527 249 568 252
rect 572 249 613 252
rect 617 249 658 252
rect 662 249 703 252
rect 707 249 748 252
rect 752 249 793 252
rect 797 249 838 252
rect 842 249 883 252
rect 887 249 900 252
rect 0 232 34 235
rect 38 232 79 235
rect 83 232 124 235
rect 128 232 169 235
rect 173 232 214 235
rect 218 232 259 235
rect 263 232 304 235
rect 308 232 349 235
rect 353 232 394 235
rect 398 232 439 235
rect 443 232 484 235
rect 488 232 529 235
rect 533 232 574 235
rect 578 232 619 235
rect 623 232 664 235
rect 668 232 709 235
rect 713 232 754 235
rect 758 232 799 235
rect 803 232 844 235
rect 848 232 889 235
rect 893 232 900 235
rect 0 225 19 228
rect 23 225 64 228
rect 68 225 109 228
rect 113 225 154 228
rect 158 225 199 228
rect 203 225 244 228
rect 248 225 289 228
rect 293 225 334 228
rect 338 225 379 228
rect 383 225 424 228
rect 428 225 469 228
rect 473 225 514 228
rect 518 225 559 228
rect 563 225 604 228
rect 608 225 649 228
rect 653 225 694 228
rect 698 225 739 228
rect 743 225 784 228
rect 788 225 829 228
rect 833 225 874 228
rect 878 225 900 228
rect 0 204 28 207
rect 32 204 73 207
rect 77 204 118 207
rect 122 204 163 207
rect 167 204 208 207
rect 212 204 253 207
rect 257 204 298 207
rect 302 204 343 207
rect 347 204 388 207
rect 392 204 433 207
rect 437 204 478 207
rect 482 204 523 207
rect 527 204 568 207
rect 572 204 613 207
rect 617 204 658 207
rect 662 204 703 207
rect 707 204 748 207
rect 752 204 793 207
rect 797 204 838 207
rect 842 204 883 207
rect 887 204 900 207
rect 0 187 34 190
rect 38 187 79 190
rect 83 187 124 190
rect 128 187 169 190
rect 173 187 214 190
rect 218 187 259 190
rect 263 187 304 190
rect 308 187 349 190
rect 353 187 394 190
rect 398 187 439 190
rect 443 187 484 190
rect 488 187 529 190
rect 533 187 574 190
rect 578 187 619 190
rect 623 187 664 190
rect 668 187 709 190
rect 713 187 754 190
rect 758 187 799 190
rect 803 187 844 190
rect 848 187 889 190
rect 893 187 900 190
rect 0 180 19 183
rect 23 180 64 183
rect 68 180 109 183
rect 113 180 154 183
rect 158 180 199 183
rect 203 180 244 183
rect 248 180 289 183
rect 293 180 334 183
rect 338 180 379 183
rect 383 180 424 183
rect 428 180 469 183
rect 473 180 514 183
rect 518 180 559 183
rect 563 180 604 183
rect 608 180 649 183
rect 653 180 694 183
rect 698 180 739 183
rect 743 180 784 183
rect 788 180 829 183
rect 833 180 874 183
rect 878 180 900 183
rect 0 159 28 162
rect 32 159 73 162
rect 77 159 118 162
rect 122 159 163 162
rect 167 159 208 162
rect 212 159 253 162
rect 257 159 298 162
rect 302 159 343 162
rect 347 159 388 162
rect 392 159 433 162
rect 437 159 478 162
rect 482 159 523 162
rect 527 159 568 162
rect 572 159 613 162
rect 617 159 658 162
rect 662 159 703 162
rect 707 159 748 162
rect 752 159 793 162
rect 797 159 838 162
rect 842 159 883 162
rect 887 159 900 162
rect 0 142 34 145
rect 38 142 79 145
rect 83 142 124 145
rect 128 142 169 145
rect 173 142 214 145
rect 218 142 259 145
rect 263 142 304 145
rect 308 142 349 145
rect 353 142 394 145
rect 398 142 439 145
rect 443 142 484 145
rect 488 142 529 145
rect 533 142 574 145
rect 578 142 619 145
rect 623 142 664 145
rect 668 142 709 145
rect 713 142 754 145
rect 758 142 799 145
rect 803 142 844 145
rect 848 142 889 145
rect 893 142 900 145
rect 0 135 19 138
rect 23 135 64 138
rect 68 135 109 138
rect 113 135 154 138
rect 158 135 199 138
rect 203 135 244 138
rect 248 135 289 138
rect 293 135 334 138
rect 338 135 379 138
rect 383 135 424 138
rect 428 135 469 138
rect 473 135 514 138
rect 518 135 559 138
rect 563 135 604 138
rect 608 135 649 138
rect 653 135 694 138
rect 698 135 739 138
rect 743 135 784 138
rect 788 135 829 138
rect 833 135 874 138
rect 878 135 900 138
rect 0 114 28 117
rect 32 114 73 117
rect 77 114 118 117
rect 122 114 163 117
rect 167 114 208 117
rect 212 114 253 117
rect 257 114 298 117
rect 302 114 343 117
rect 347 114 388 117
rect 392 114 433 117
rect 437 114 478 117
rect 482 114 523 117
rect 527 114 568 117
rect 572 114 613 117
rect 617 114 658 117
rect 662 114 703 117
rect 707 114 748 117
rect 752 114 793 117
rect 797 114 838 117
rect 842 114 883 117
rect 887 114 900 117
rect 0 97 34 100
rect 38 97 79 100
rect 83 97 124 100
rect 128 97 169 100
rect 173 97 214 100
rect 218 97 259 100
rect 263 97 304 100
rect 308 97 349 100
rect 353 97 394 100
rect 398 97 439 100
rect 443 97 484 100
rect 488 97 529 100
rect 533 97 574 100
rect 578 97 619 100
rect 623 97 664 100
rect 668 97 709 100
rect 713 97 754 100
rect 758 97 799 100
rect 803 97 844 100
rect 848 97 889 100
rect 893 97 900 100
rect 0 90 19 93
rect 23 90 64 93
rect 68 90 109 93
rect 113 90 154 93
rect 158 90 199 93
rect 203 90 244 93
rect 248 90 289 93
rect 293 90 334 93
rect 338 90 379 93
rect 383 90 424 93
rect 428 90 469 93
rect 473 90 514 93
rect 518 90 559 93
rect 563 90 604 93
rect 608 90 649 93
rect 653 90 694 93
rect 698 90 739 93
rect 743 90 784 93
rect 788 90 829 93
rect 833 90 874 93
rect 878 90 900 93
rect 0 69 28 72
rect 32 69 73 72
rect 77 69 118 72
rect 122 69 163 72
rect 167 69 208 72
rect 212 69 253 72
rect 257 69 298 72
rect 302 69 343 72
rect 347 69 388 72
rect 392 69 433 72
rect 437 69 478 72
rect 482 69 523 72
rect 527 69 568 72
rect 572 69 613 72
rect 617 69 658 72
rect 662 69 703 72
rect 707 69 748 72
rect 752 69 793 72
rect 797 69 838 72
rect 842 69 883 72
rect 887 69 900 72
rect 0 52 34 55
rect 38 52 79 55
rect 83 52 124 55
rect 128 52 169 55
rect 173 52 214 55
rect 218 52 259 55
rect 263 52 304 55
rect 308 52 349 55
rect 353 52 394 55
rect 398 52 439 55
rect 443 52 484 55
rect 488 52 529 55
rect 533 52 574 55
rect 578 52 619 55
rect 623 52 664 55
rect 668 52 709 55
rect 713 52 754 55
rect 758 52 799 55
rect 803 52 844 55
rect 848 52 889 55
rect 893 52 900 55
rect 0 45 19 48
rect 23 45 64 48
rect 68 45 109 48
rect 113 45 154 48
rect 158 45 199 48
rect 203 45 244 48
rect 248 45 289 48
rect 293 45 334 48
rect 338 45 379 48
rect 383 45 424 48
rect 428 45 469 48
rect 473 45 514 48
rect 518 45 559 48
rect 563 45 604 48
rect 608 45 649 48
rect 653 45 694 48
rect 698 45 739 48
rect 743 45 784 48
rect 788 45 829 48
rect 833 45 874 48
rect 878 45 900 48
rect 0 24 28 27
rect 32 24 73 27
rect 77 24 118 27
rect 122 24 163 27
rect 167 24 208 27
rect 212 24 253 27
rect 257 24 298 27
rect 302 24 343 27
rect 347 24 388 27
rect 392 24 433 27
rect 437 24 478 27
rect 482 24 523 27
rect 527 24 568 27
rect 572 24 613 27
rect 617 24 658 27
rect 662 24 703 27
rect 707 24 748 27
rect 752 24 793 27
rect 797 24 838 27
rect 842 24 883 27
rect 887 24 900 27
rect 0 7 34 10
rect 38 7 79 10
rect 83 7 124 10
rect 128 7 169 10
rect 173 7 214 10
rect 218 7 259 10
rect 263 7 304 10
rect 308 7 349 10
rect 353 7 394 10
rect 398 7 439 10
rect 443 7 484 10
rect 488 7 529 10
rect 533 7 574 10
rect 578 7 619 10
rect 623 7 664 10
rect 668 7 709 10
rect 713 7 754 10
rect 758 7 799 10
rect 803 7 844 10
rect 848 7 889 10
rect 893 7 900 10
rect 0 0 19 3
rect 23 0 64 3
rect 68 0 109 3
rect 113 0 154 3
rect 158 0 199 3
rect 203 0 244 3
rect 248 0 289 3
rect 293 0 334 3
rect 338 0 379 3
rect 383 0 424 3
rect 428 0 469 3
rect 473 0 514 3
rect 518 0 559 3
rect 563 0 604 3
rect 608 0 649 3
rect 653 0 694 3
rect 698 0 739 3
rect 743 0 784 3
rect 788 0 829 3
rect 833 0 874 3
rect 878 0 900 3
rect -216 -157 -188 -154
rect -304 -161 -300 -157
rect -184 -157 -171 -154
rect -280 -169 -277 -165
rect -216 -174 -182 -171
rect -178 -174 -171 -171
rect -268 -179 -257 -175
rect -216 -181 -197 -178
rect -193 -181 -171 -178
<< metal3 >>
rect -306 -151 -271 -116
<< end >>
