magic
tech scmos
timestamp 1354245769
use pixel_2.1  pixel_2.1_0
array 0 31 96 0 31 96
timestamp 1354245571
transform 1 0 0 0 1 0
box 0 0 96 96
<< end >>
