magic
tech scmos
timestamp 1355258800
<< nwell >>
rect -20 86 152 121
<< pwell >>
rect -1 51 133 86
<< ntransistor >>
rect 25 57 29 77
rect 35 57 39 77
rect 45 57 49 77
rect 55 57 59 77
rect 73 57 77 77
rect 83 57 87 77
rect 93 57 97 77
rect 103 57 107 77
<< ptransistor >>
rect -3 95 1 115
rect 7 95 11 115
rect 25 95 29 115
rect 35 95 39 115
rect 45 95 49 115
rect 55 95 59 115
rect 73 95 77 115
rect 83 95 87 115
rect 93 95 97 115
rect 103 95 107 115
rect 121 95 125 115
rect 131 95 135 115
<< ndiffusion >>
rect 24 57 25 77
rect 29 57 30 77
rect 34 57 35 77
rect 39 57 40 77
rect 44 57 45 77
rect 49 57 50 77
rect 54 57 55 77
rect 59 57 60 77
rect 72 57 73 77
rect 77 57 78 77
rect 82 57 83 77
rect 87 57 88 77
rect 92 57 93 77
rect 97 57 98 77
rect 102 57 103 77
rect 107 57 108 77
<< pdiffusion >>
rect -10 95 -8 115
rect -4 95 -3 115
rect 1 95 2 115
rect 6 95 7 115
rect 11 95 12 115
rect 24 95 25 115
rect 29 95 30 115
rect 34 95 35 115
rect 39 95 40 115
rect 44 95 45 115
rect 49 95 50 115
rect 54 95 55 115
rect 59 95 60 115
rect 72 95 73 115
rect 77 95 78 115
rect 82 95 83 115
rect 87 95 88 115
rect 92 95 93 115
rect 97 95 98 115
rect 102 95 103 115
rect 107 95 108 115
rect 120 95 121 115
rect 125 95 126 115
rect 130 95 131 115
rect 135 95 136 115
rect 140 95 142 115
<< ndcontact >>
rect 20 57 24 77
rect 30 57 34 77
rect 40 57 44 77
rect 50 57 54 77
rect 60 57 64 77
rect 68 57 72 77
rect 78 57 82 77
rect 88 57 92 77
rect 98 57 102 77
rect 108 57 112 77
<< pdcontact >>
rect -8 95 -4 115
rect 2 95 6 115
rect 12 95 16 115
rect 20 95 24 115
rect 30 95 34 115
rect 40 95 44 115
rect 50 95 54 115
rect 60 95 64 115
rect 68 95 72 115
rect 78 95 82 115
rect 88 95 92 115
rect 98 95 102 115
rect 108 95 112 115
rect 116 95 120 115
rect 126 95 130 115
rect 136 95 140 115
<< psubstratepdiff >>
rect 3 76 20 77
rect 3 58 5 76
rect 19 58 20 76
rect 3 57 20 58
rect 112 76 129 77
rect 112 58 113 76
rect 127 58 129 76
rect 112 57 129 58
<< nsubstratendiff >>
rect -11 95 -10 115
rect 142 95 143 115
<< psubstratepcontact >>
rect 5 58 19 76
rect 113 58 127 76
<< nsubstratencontact >>
rect -15 95 -11 115
rect 143 95 147 115
<< polysilicon >>
rect 9 121 123 123
rect 9 118 11 121
rect -20 116 11 118
rect 121 118 123 121
rect -3 115 1 116
rect 7 115 11 116
rect 25 115 29 117
rect 35 115 39 117
rect 45 115 49 117
rect 55 115 59 117
rect 73 115 77 117
rect 83 115 87 117
rect 93 115 97 117
rect 103 115 107 117
rect 121 116 152 118
rect 121 115 125 116
rect 131 115 135 116
rect -3 93 1 95
rect 7 93 11 95
rect 25 94 29 95
rect 35 94 39 95
rect 25 92 39 94
rect 45 94 49 95
rect 55 94 59 95
rect 45 93 59 94
rect 45 92 53 93
rect 37 89 39 92
rect 57 92 59 93
rect 73 94 77 95
rect 83 94 87 95
rect 73 93 87 94
rect 73 92 75 93
rect 79 92 87 93
rect 93 94 97 95
rect 103 94 107 95
rect 93 92 107 94
rect 121 93 125 95
rect 131 93 135 95
rect 93 89 95 92
rect -20 87 39 89
rect 37 85 39 87
rect 93 87 152 89
rect 93 85 95 87
rect 37 83 95 85
rect 25 79 27 83
rect 105 79 107 83
rect 25 77 29 79
rect 35 77 39 79
rect 45 77 49 79
rect 55 77 59 79
rect 73 77 77 79
rect 83 77 87 79
rect 93 77 97 79
rect 103 77 107 79
rect 25 56 29 57
rect 35 56 39 57
rect 45 56 49 57
rect 55 56 59 57
rect 25 54 59 56
rect 73 56 77 57
rect 83 56 87 57
rect 93 56 97 57
rect 103 56 107 57
rect 73 54 107 56
<< polycontact >>
rect 53 89 57 93
rect 75 89 79 93
rect 27 79 31 83
rect 101 79 105 83
<< metal1 >>
rect 12 125 120 128
rect 12 121 16 125
rect 116 121 120 125
rect -8 118 16 121
rect -8 115 -4 118
rect 12 115 16 118
rect -11 95 -8 115
rect 20 118 64 121
rect 20 115 24 118
rect 40 115 44 118
rect 60 115 64 118
rect 2 92 6 95
rect 20 92 24 95
rect 2 89 24 92
rect 68 118 112 121
rect 68 115 72 118
rect 88 115 92 118
rect 108 115 112 118
rect 30 83 34 95
rect 31 79 34 83
rect 30 77 34 79
rect 50 93 54 95
rect 78 93 82 95
rect 50 89 53 93
rect 50 86 64 89
rect 79 89 82 93
rect 68 86 82 89
rect 50 77 54 86
rect 78 77 82 86
rect 98 83 102 95
rect 116 118 140 121
rect 116 115 120 118
rect 136 115 140 118
rect 140 95 143 115
rect 108 92 112 95
rect 126 92 130 95
rect 108 89 130 92
rect 98 79 101 83
rect 98 77 102 79
rect 19 58 20 76
rect 20 54 24 57
rect 40 54 44 57
rect 60 54 64 57
rect 112 58 113 76
rect 68 54 72 57
rect 88 54 92 57
rect 108 54 112 57
rect 20 51 112 54
<< m2contact >>
rect -20 95 -15 115
rect 64 86 68 90
rect 147 95 152 115
rect 1 58 5 76
rect 127 58 131 76
<< metal2 >>
rect 64 90 68 128
rect -20 58 1 76
rect 131 58 152 76
<< end >>
