magic
tech scmos
timestamp 1355359077
<< nsubstratencontact >>
rect 663 688 667 692
<< metal1 >>
rect 629 4481 669 4491
rect 662 4275 669 4481
rect 662 4260 4217 4275
<< metal2 >>
rect 649 4259 652 4269
rect 655 4259 658 4269
rect 4332 625 4336 635
rect 4243 594 4248 614
rect 4420 594 4425 614
<< m3contact >>
rect 596 4466 612 4487
rect 606 571 633 589
<< metal3 >>
rect 543 4487 658 4488
rect 543 4466 596 4487
rect 612 4466 658 4487
rect 543 702 658 4466
rect 543 589 4220 702
rect 543 571 606 589
rect 633 576 4220 589
rect 633 571 4420 576
rect 543 556 4420 571
rect 543 550 4220 556
use blankpad  blankpad_11
timestamp 1259953556
transform -1 0 841 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_12
timestamp 1259953556
transform -1 0 1315 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_13
timestamp 1259953556
transform -1 0 1789 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_14
timestamp 1259953556
transform -1 0 2263 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_15
timestamp 1259953556
transform -1 0 2737 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_16
timestamp 1259953556
transform -1 0 3211 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_17
timestamp 1259953556
transform -1 0 3685 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_10
timestamp 1259953556
transform -1 0 4159 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_9
timestamp 1259953556
transform -1 0 4633 0 -1 5000
box -2 0 476 513
use padframe_top  padframe_top_0
timestamp 1259953556
transform 1 0 0 0 1 4487
box 0 0 5000 513
use blankpad  blankpad_27
timestamp 1259953556
transform 0 1 0 -1 0 4633
box -2 0 476 513
use blankpad  blankpad_28
timestamp 1259953556
transform 0 1 0 -1 0 4159
box -2 0 476 513
use blankpad  blankpad_35
timestamp 1259953556
transform 0 1 0 -1 0 3685
box -2 0 476 513
use blankpad  blankpad_34
timestamp 1259953556
transform 0 1 0 -1 0 3211
box -2 0 476 513
use blankpad  blankpad_33
timestamp 1259953556
transform 0 1 0 -1 0 2737
box -2 0 476 513
use blankpad  blankpad_32
timestamp 1259953556
transform 0 1 0 -1 0 2263
box -2 0 476 513
use blankpad  blankpad_31
timestamp 1259953556
transform 0 1 0 -1 0 1789
box -2 0 476 513
use blankpad  blankpad_30
timestamp 1259953556
transform 0 1 0 -1 0 1315
box -2 0 476 513
use imager_nopads  imager_nopads_0
timestamp 1355359077
transform 1 0 662 0 1 705
box -116 -152 3558 3579
use blankpad  blankpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 4159
box -2 0 476 513
use blankpad  blankpad_3
timestamp 1259953556
transform 0 -1 5000 1 0 3685
box -2 0 476 513
use blankpad  blankpad_4
timestamp 1259953556
transform 0 -1 5000 1 0 3211
box -2 0 476 513
use blankpad  blankpad_5
timestamp 1259953556
transform 0 -1 5000 1 0 2737
box -2 0 476 513
use blankpad  blankpad_6
timestamp 1259953556
transform 0 -1 5000 1 0 2263
box -2 0 476 513
use blankpad  blankpad_7
timestamp 1259953556
transform 0 -1 5000 1 0 1789
box -2 0 476 513
use blankpad  blankpad_8
timestamp 1259953556
transform 0 -1 5000 1 0 1315
box -2 0 476 513
use blankpad  blankpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 841
box -2 0 476 513
use diffamp  diffamp_0
timestamp 1355272872
transform 1 0 4268 0 1 499
box -20 51 152 128
use padframe_left  padframe_left_0
timestamp 1259953556
transform 1 0 0 0 1 367
box 2 2 513 4264
use blankpad  blankpad_29
timestamp 1259953556
transform 0 1 0 -1 0 841
box -2 0 476 513
use blankpad  blankpad_18
timestamp 1259953556
transform 1 0 367 0 1 0
box -2 0 476 513
use blankpad  blankpad_19
timestamp 1259953556
transform 1 0 841 0 1 0
box -2 0 476 513
use blankpad  blankpad_26
timestamp 1259953556
transform 1 0 1315 0 1 0
box -2 0 476 513
use blankpad  blankpad_25
timestamp 1259953556
transform 1 0 1789 0 1 0
box -2 0 476 513
use blankpad  blankpad_24
timestamp 1259953556
transform 1 0 2263 0 1 0
box -2 0 476 513
use blankpad  blankpad_23
timestamp 1259953556
transform 1 0 2737 0 1 0
box -2 0 476 513
use blankpad  blankpad_22
timestamp 1259953556
transform 1 0 3211 0 1 0
box -2 0 476 513
use blankpad  blankpad_21
timestamp 1259953556
transform 1 0 3685 0 1 0
box -2 0 476 513
use padframe_right  padframe_right_0
timestamp 1259953556
transform 1 0 4487 0 1 367
box 0 2 511 4264
use blankpad  blankpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 367
box -2 0 476 513
use blankpad  blankpad_20
timestamp 1259953556
transform 1 0 4159 0 1 0
box -2 0 476 513
use padframe_bottom  padframe_bottom_0
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 5000 513
<< end >>
