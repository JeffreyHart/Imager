magic
tech scmos
timestamp 1354597133
use csrlend  csrlend_0
timestamp 1348671188
transform 1 0 -25 0 1 -152
box 0 11 20 81
use csrldff  csrldff_0
array 0 63 48 0 0 96
timestamp 1354594767
transform 1 0 8 0 1 -152
box -13 0 35 96
<< end >>
