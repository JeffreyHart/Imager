magic
tech scmos
timestamp 1354596218
<< nwell >>
rect -3 -23 25 -6
rect 74 -23 121 -6
rect 170 -23 217 -6
rect 266 -23 313 -6
rect 362 -23 409 -6
rect 458 -23 505 -6
rect 554 -23 601 -6
rect 650 -23 697 -6
rect 746 -23 793 -6
rect 842 -23 889 -6
rect 938 -23 966 -6
<< pwell >>
rect -3 -6 966 99
rect 25 -23 74 -6
rect 121 -23 170 -6
rect 217 -23 266 -6
rect 313 -23 362 -6
rect 409 -23 458 -6
rect 505 -23 554 -6
rect 601 -23 650 -6
rect 697 -23 746 -6
rect 793 -23 842 -6
rect 889 -23 938 -6
rect -3 -56 966 -23
<< ntransistor >>
rect 27 66 30 68
rect 14 59 16 62
rect 69 66 72 68
rect 53 59 56 60
rect 83 59 85 62
rect 23 50 25 53
rect 33 50 35 53
rect 64 50 66 53
rect 74 50 76 53
rect 123 66 126 68
rect 110 59 112 62
rect 165 66 168 68
rect 149 59 152 60
rect 179 59 181 62
rect 119 50 121 53
rect 129 50 131 53
rect 23 40 25 43
rect 33 40 35 43
rect 160 50 162 53
rect 170 50 172 53
rect 219 66 222 68
rect 206 59 208 62
rect 261 66 264 68
rect 245 59 248 60
rect 275 59 277 62
rect 215 50 217 53
rect 225 50 227 53
rect 64 40 66 43
rect 74 40 76 43
rect 14 31 16 34
rect 53 33 56 34
rect 27 25 30 27
rect 83 31 85 34
rect 69 25 72 27
rect 119 40 121 43
rect 129 40 131 43
rect 256 50 258 53
rect 266 50 268 53
rect 315 66 318 68
rect 302 59 304 62
rect 357 66 360 68
rect 341 59 344 60
rect 371 59 373 62
rect 311 50 313 53
rect 321 50 323 53
rect 160 40 162 43
rect 170 40 172 43
rect 110 31 112 34
rect 149 33 152 34
rect 123 25 126 27
rect 179 31 181 34
rect 165 25 168 27
rect 215 40 217 43
rect 225 40 227 43
rect 352 50 354 53
rect 362 50 364 53
rect 411 66 414 68
rect 398 59 400 62
rect 453 66 456 68
rect 437 59 440 60
rect 467 59 469 62
rect 407 50 409 53
rect 417 50 419 53
rect 256 40 258 43
rect 266 40 268 43
rect 206 31 208 34
rect 245 33 248 34
rect 219 25 222 27
rect 275 31 277 34
rect 261 25 264 27
rect 311 40 313 43
rect 321 40 323 43
rect 448 50 450 53
rect 458 50 460 53
rect 507 66 510 68
rect 494 59 496 62
rect 549 66 552 68
rect 533 59 536 60
rect 563 59 565 62
rect 503 50 505 53
rect 513 50 515 53
rect 352 40 354 43
rect 362 40 364 43
rect 302 31 304 34
rect 341 33 344 34
rect 315 25 318 27
rect 371 31 373 34
rect 357 25 360 27
rect 407 40 409 43
rect 417 40 419 43
rect 544 50 546 53
rect 554 50 556 53
rect 603 66 606 68
rect 590 59 592 62
rect 645 66 648 68
rect 629 59 632 60
rect 659 59 661 62
rect 599 50 601 53
rect 609 50 611 53
rect 448 40 450 43
rect 458 40 460 43
rect 398 31 400 34
rect 437 33 440 34
rect 411 25 414 27
rect 467 31 469 34
rect 453 25 456 27
rect 503 40 505 43
rect 513 40 515 43
rect 640 50 642 53
rect 650 50 652 53
rect 699 66 702 68
rect 686 59 688 62
rect 741 66 744 68
rect 725 59 728 60
rect 755 59 757 62
rect 695 50 697 53
rect 705 50 707 53
rect 544 40 546 43
rect 554 40 556 43
rect 494 31 496 34
rect 533 33 536 34
rect 507 25 510 27
rect 563 31 565 34
rect 549 25 552 27
rect 599 40 601 43
rect 609 40 611 43
rect 736 50 738 53
rect 746 50 748 53
rect 795 66 798 68
rect 782 59 784 62
rect 837 66 840 68
rect 821 59 824 60
rect 851 59 853 62
rect 791 50 793 53
rect 801 50 803 53
rect 640 40 642 43
rect 650 40 652 43
rect 590 31 592 34
rect 629 33 632 34
rect 603 25 606 27
rect 659 31 661 34
rect 645 25 648 27
rect 695 40 697 43
rect 705 40 707 43
rect 832 50 834 53
rect 842 50 844 53
rect 891 66 894 68
rect 878 59 880 62
rect 933 66 936 68
rect 917 59 920 60
rect 947 59 949 62
rect 887 50 889 53
rect 897 50 899 53
rect 736 40 738 43
rect 746 40 748 43
rect 686 31 688 34
rect 725 33 728 34
rect 699 25 702 27
rect 755 31 757 34
rect 741 25 744 27
rect 791 40 793 43
rect 801 40 803 43
rect 928 50 930 53
rect 938 50 940 53
rect 832 40 834 43
rect 842 40 844 43
rect 782 31 784 34
rect 821 33 824 34
rect 795 25 798 27
rect 851 31 853 34
rect 837 25 840 27
rect 887 40 889 43
rect 897 40 899 43
rect 928 40 930 43
rect 938 40 940 43
rect 878 31 880 34
rect 917 33 920 34
rect 891 25 894 27
rect 947 31 949 34
rect 933 25 936 27
rect 37 -16 39 -13
rect 60 -16 62 -13
rect 133 -16 135 -13
rect 29 -32 31 -29
rect 9 -40 11 -37
rect 14 -40 16 -37
rect 37 -32 39 -29
rect 156 -16 158 -13
rect 229 -16 231 -13
rect 60 -32 62 -29
rect 68 -32 70 -29
rect 125 -32 127 -29
rect 83 -40 85 -37
rect 88 -40 90 -37
rect 105 -40 107 -37
rect 110 -40 112 -37
rect 133 -32 135 -29
rect 252 -16 254 -13
rect 325 -16 327 -13
rect 156 -32 158 -29
rect 164 -32 166 -29
rect 221 -32 223 -29
rect 179 -40 181 -37
rect 184 -40 186 -37
rect 201 -40 203 -37
rect 206 -40 208 -37
rect 229 -32 231 -29
rect 348 -16 350 -13
rect 421 -16 423 -13
rect 252 -32 254 -29
rect 260 -32 262 -29
rect 317 -32 319 -29
rect 275 -40 277 -37
rect 280 -40 282 -37
rect 297 -40 299 -37
rect 302 -40 304 -37
rect 325 -32 327 -29
rect 444 -16 446 -13
rect 517 -16 519 -13
rect 348 -32 350 -29
rect 356 -32 358 -29
rect 413 -32 415 -29
rect 371 -40 373 -37
rect 376 -40 378 -37
rect 393 -40 395 -37
rect 398 -40 400 -37
rect 421 -32 423 -29
rect 540 -16 542 -13
rect 613 -16 615 -13
rect 444 -32 446 -29
rect 452 -32 454 -29
rect 509 -32 511 -29
rect 467 -40 469 -37
rect 472 -40 474 -37
rect 489 -40 491 -37
rect 494 -40 496 -37
rect 517 -32 519 -29
rect 636 -16 638 -13
rect 709 -16 711 -13
rect 540 -32 542 -29
rect 548 -32 550 -29
rect 605 -32 607 -29
rect 563 -40 565 -37
rect 568 -40 570 -37
rect 585 -40 587 -37
rect 590 -40 592 -37
rect 613 -32 615 -29
rect 732 -16 734 -13
rect 805 -16 807 -13
rect 636 -32 638 -29
rect 644 -32 646 -29
rect 701 -32 703 -29
rect 659 -40 661 -37
rect 664 -40 666 -37
rect 681 -40 683 -37
rect 686 -40 688 -37
rect 709 -32 711 -29
rect 828 -16 830 -13
rect 901 -16 903 -13
rect 732 -32 734 -29
rect 740 -32 742 -29
rect 797 -32 799 -29
rect 755 -40 757 -37
rect 760 -40 762 -37
rect 777 -40 779 -37
rect 782 -40 784 -37
rect 805 -32 807 -29
rect 924 -16 926 -13
rect 828 -32 830 -29
rect 836 -32 838 -29
rect 893 -32 895 -29
rect 851 -40 853 -37
rect 856 -40 858 -37
rect 873 -40 875 -37
rect 878 -40 880 -37
rect 901 -32 903 -29
rect 924 -32 926 -29
rect 932 -32 934 -29
rect 947 -40 949 -37
rect 952 -40 954 -37
<< ptransistor >>
rect 12 -16 14 -13
rect 85 -16 87 -13
rect 108 -16 110 -13
rect 181 -16 183 -13
rect 204 -16 206 -13
rect 277 -16 279 -13
rect 300 -16 302 -13
rect 373 -16 375 -13
rect 396 -16 398 -13
rect 469 -16 471 -13
rect 492 -16 494 -13
rect 565 -16 567 -13
rect 588 -16 590 -13
rect 661 -16 663 -13
rect 684 -16 686 -13
rect 757 -16 759 -13
rect 780 -16 782 -13
rect 853 -16 855 -13
rect 876 -16 878 -13
rect 949 -16 951 -13
<< ndiffusion >>
rect 3 70 48 93
rect 3 66 19 70
rect 25 69 48 70
rect 3 62 13 66
rect 27 68 30 69
rect 27 65 30 66
rect 3 59 14 62
rect 16 59 17 62
rect 3 57 12 59
rect 3 51 9 57
rect 35 61 48 69
rect 51 70 96 93
rect 51 69 74 70
rect 51 61 64 69
rect 69 68 72 69
rect 69 65 72 66
rect 80 66 96 70
rect 86 62 96 66
rect 35 59 46 61
rect 53 60 64 61
rect 56 59 64 60
rect 82 59 83 62
rect 85 59 96 62
rect 87 57 96 59
rect 3 48 13 51
rect 21 50 23 53
rect 25 50 33 53
rect 35 50 36 53
rect 63 50 64 53
rect 66 50 74 53
rect 76 50 78 53
rect 90 51 96 57
rect 86 48 96 51
rect 99 70 144 93
rect 99 66 115 70
rect 121 69 144 70
rect 99 62 109 66
rect 123 68 126 69
rect 123 65 126 66
rect 99 59 110 62
rect 112 59 113 62
rect 99 57 108 59
rect 99 51 105 57
rect 131 61 144 69
rect 147 70 192 93
rect 147 69 170 70
rect 147 61 160 69
rect 165 68 168 69
rect 165 65 168 66
rect 176 66 192 70
rect 182 62 192 66
rect 131 59 142 61
rect 149 60 160 61
rect 152 59 160 60
rect 178 59 179 62
rect 181 59 192 62
rect 183 57 192 59
rect 99 48 109 51
rect 117 50 119 53
rect 121 50 129 53
rect 131 50 132 53
rect 3 42 13 45
rect 3 36 9 42
rect 21 40 23 43
rect 25 40 33 43
rect 35 40 36 43
rect 3 34 12 36
rect 159 50 160 53
rect 162 50 170 53
rect 172 50 174 53
rect 186 51 192 57
rect 182 48 192 51
rect 195 70 240 93
rect 195 66 211 70
rect 217 69 240 70
rect 195 62 205 66
rect 219 68 222 69
rect 219 65 222 66
rect 195 59 206 62
rect 208 59 209 62
rect 195 57 204 59
rect 195 51 201 57
rect 227 61 240 69
rect 243 70 288 93
rect 243 69 266 70
rect 243 61 256 69
rect 261 68 264 69
rect 261 65 264 66
rect 272 66 288 70
rect 278 62 288 66
rect 227 59 238 61
rect 245 60 256 61
rect 248 59 256 60
rect 274 59 275 62
rect 277 59 288 62
rect 279 57 288 59
rect 195 48 205 51
rect 213 50 215 53
rect 217 50 225 53
rect 227 50 228 53
rect 63 40 64 43
rect 66 40 74 43
rect 76 40 78 43
rect 86 42 96 45
rect 3 31 14 34
rect 16 31 17 34
rect 35 32 46 34
rect 56 33 64 34
rect 53 32 64 33
rect 3 27 13 31
rect 3 23 19 27
rect 27 27 30 28
rect 27 24 30 25
rect 35 24 48 32
rect 25 23 48 24
rect 3 0 48 23
rect 51 24 64 32
rect 90 36 96 42
rect 87 34 96 36
rect 82 31 83 34
rect 85 31 96 34
rect 69 27 72 28
rect 69 24 72 25
rect 86 27 96 31
rect 51 23 74 24
rect 80 23 96 27
rect 51 0 96 23
rect 99 42 109 45
rect 99 36 105 42
rect 117 40 119 43
rect 121 40 129 43
rect 131 40 132 43
rect 99 34 108 36
rect 255 50 256 53
rect 258 50 266 53
rect 268 50 270 53
rect 282 51 288 57
rect 278 48 288 51
rect 291 70 336 93
rect 291 66 307 70
rect 313 69 336 70
rect 291 62 301 66
rect 315 68 318 69
rect 315 65 318 66
rect 291 59 302 62
rect 304 59 305 62
rect 291 57 300 59
rect 291 51 297 57
rect 323 61 336 69
rect 339 70 384 93
rect 339 69 362 70
rect 339 61 352 69
rect 357 68 360 69
rect 357 65 360 66
rect 368 66 384 70
rect 374 62 384 66
rect 323 59 334 61
rect 341 60 352 61
rect 344 59 352 60
rect 370 59 371 62
rect 373 59 384 62
rect 375 57 384 59
rect 291 48 301 51
rect 309 50 311 53
rect 313 50 321 53
rect 323 50 324 53
rect 159 40 160 43
rect 162 40 170 43
rect 172 40 174 43
rect 182 42 192 45
rect 99 31 110 34
rect 112 31 113 34
rect 131 32 142 34
rect 152 33 160 34
rect 149 32 160 33
rect 99 27 109 31
rect 99 23 115 27
rect 123 27 126 28
rect 123 24 126 25
rect 131 24 144 32
rect 121 23 144 24
rect 99 0 144 23
rect 147 24 160 32
rect 186 36 192 42
rect 183 34 192 36
rect 178 31 179 34
rect 181 31 192 34
rect 165 27 168 28
rect 165 24 168 25
rect 182 27 192 31
rect 147 23 170 24
rect 176 23 192 27
rect 147 0 192 23
rect 195 42 205 45
rect 195 36 201 42
rect 213 40 215 43
rect 217 40 225 43
rect 227 40 228 43
rect 195 34 204 36
rect 351 50 352 53
rect 354 50 362 53
rect 364 50 366 53
rect 378 51 384 57
rect 374 48 384 51
rect 387 70 432 93
rect 387 66 403 70
rect 409 69 432 70
rect 387 62 397 66
rect 411 68 414 69
rect 411 65 414 66
rect 387 59 398 62
rect 400 59 401 62
rect 387 57 396 59
rect 387 51 393 57
rect 419 61 432 69
rect 435 70 480 93
rect 435 69 458 70
rect 435 61 448 69
rect 453 68 456 69
rect 453 65 456 66
rect 464 66 480 70
rect 470 62 480 66
rect 419 59 430 61
rect 437 60 448 61
rect 440 59 448 60
rect 466 59 467 62
rect 469 59 480 62
rect 471 57 480 59
rect 387 48 397 51
rect 405 50 407 53
rect 409 50 417 53
rect 419 50 420 53
rect 255 40 256 43
rect 258 40 266 43
rect 268 40 270 43
rect 278 42 288 45
rect 195 31 206 34
rect 208 31 209 34
rect 227 32 238 34
rect 248 33 256 34
rect 245 32 256 33
rect 195 27 205 31
rect 195 23 211 27
rect 219 27 222 28
rect 219 24 222 25
rect 227 24 240 32
rect 217 23 240 24
rect 195 0 240 23
rect 243 24 256 32
rect 282 36 288 42
rect 279 34 288 36
rect 274 31 275 34
rect 277 31 288 34
rect 261 27 264 28
rect 261 24 264 25
rect 278 27 288 31
rect 243 23 266 24
rect 272 23 288 27
rect 243 0 288 23
rect 291 42 301 45
rect 291 36 297 42
rect 309 40 311 43
rect 313 40 321 43
rect 323 40 324 43
rect 291 34 300 36
rect 447 50 448 53
rect 450 50 458 53
rect 460 50 462 53
rect 474 51 480 57
rect 470 48 480 51
rect 483 70 528 93
rect 483 66 499 70
rect 505 69 528 70
rect 483 62 493 66
rect 507 68 510 69
rect 507 65 510 66
rect 483 59 494 62
rect 496 59 497 62
rect 483 57 492 59
rect 483 51 489 57
rect 515 61 528 69
rect 531 70 576 93
rect 531 69 554 70
rect 531 61 544 69
rect 549 68 552 69
rect 549 65 552 66
rect 560 66 576 70
rect 566 62 576 66
rect 515 59 526 61
rect 533 60 544 61
rect 536 59 544 60
rect 562 59 563 62
rect 565 59 576 62
rect 567 57 576 59
rect 483 48 493 51
rect 501 50 503 53
rect 505 50 513 53
rect 515 50 516 53
rect 351 40 352 43
rect 354 40 362 43
rect 364 40 366 43
rect 374 42 384 45
rect 291 31 302 34
rect 304 31 305 34
rect 323 32 334 34
rect 344 33 352 34
rect 341 32 352 33
rect 291 27 301 31
rect 291 23 307 27
rect 315 27 318 28
rect 315 24 318 25
rect 323 24 336 32
rect 313 23 336 24
rect 291 0 336 23
rect 339 24 352 32
rect 378 36 384 42
rect 375 34 384 36
rect 370 31 371 34
rect 373 31 384 34
rect 357 27 360 28
rect 357 24 360 25
rect 374 27 384 31
rect 339 23 362 24
rect 368 23 384 27
rect 339 0 384 23
rect 387 42 397 45
rect 387 36 393 42
rect 405 40 407 43
rect 409 40 417 43
rect 419 40 420 43
rect 387 34 396 36
rect 543 50 544 53
rect 546 50 554 53
rect 556 50 558 53
rect 570 51 576 57
rect 566 48 576 51
rect 579 70 624 93
rect 579 66 595 70
rect 601 69 624 70
rect 579 62 589 66
rect 603 68 606 69
rect 603 65 606 66
rect 579 59 590 62
rect 592 59 593 62
rect 579 57 588 59
rect 579 51 585 57
rect 611 61 624 69
rect 627 70 672 93
rect 627 69 650 70
rect 627 61 640 69
rect 645 68 648 69
rect 645 65 648 66
rect 656 66 672 70
rect 662 62 672 66
rect 611 59 622 61
rect 629 60 640 61
rect 632 59 640 60
rect 658 59 659 62
rect 661 59 672 62
rect 663 57 672 59
rect 579 48 589 51
rect 597 50 599 53
rect 601 50 609 53
rect 611 50 612 53
rect 447 40 448 43
rect 450 40 458 43
rect 460 40 462 43
rect 470 42 480 45
rect 387 31 398 34
rect 400 31 401 34
rect 419 32 430 34
rect 440 33 448 34
rect 437 32 448 33
rect 387 27 397 31
rect 387 23 403 27
rect 411 27 414 28
rect 411 24 414 25
rect 419 24 432 32
rect 409 23 432 24
rect 387 0 432 23
rect 435 24 448 32
rect 474 36 480 42
rect 471 34 480 36
rect 466 31 467 34
rect 469 31 480 34
rect 453 27 456 28
rect 453 24 456 25
rect 470 27 480 31
rect 435 23 458 24
rect 464 23 480 27
rect 435 0 480 23
rect 483 42 493 45
rect 483 36 489 42
rect 501 40 503 43
rect 505 40 513 43
rect 515 40 516 43
rect 483 34 492 36
rect 639 50 640 53
rect 642 50 650 53
rect 652 50 654 53
rect 666 51 672 57
rect 662 48 672 51
rect 675 70 720 93
rect 675 66 691 70
rect 697 69 720 70
rect 675 62 685 66
rect 699 68 702 69
rect 699 65 702 66
rect 675 59 686 62
rect 688 59 689 62
rect 675 57 684 59
rect 675 51 681 57
rect 707 61 720 69
rect 723 70 768 93
rect 723 69 746 70
rect 723 61 736 69
rect 741 68 744 69
rect 741 65 744 66
rect 752 66 768 70
rect 758 62 768 66
rect 707 59 718 61
rect 725 60 736 61
rect 728 59 736 60
rect 754 59 755 62
rect 757 59 768 62
rect 759 57 768 59
rect 675 48 685 51
rect 693 50 695 53
rect 697 50 705 53
rect 707 50 708 53
rect 543 40 544 43
rect 546 40 554 43
rect 556 40 558 43
rect 566 42 576 45
rect 483 31 494 34
rect 496 31 497 34
rect 515 32 526 34
rect 536 33 544 34
rect 533 32 544 33
rect 483 27 493 31
rect 483 23 499 27
rect 507 27 510 28
rect 507 24 510 25
rect 515 24 528 32
rect 505 23 528 24
rect 483 0 528 23
rect 531 24 544 32
rect 570 36 576 42
rect 567 34 576 36
rect 562 31 563 34
rect 565 31 576 34
rect 549 27 552 28
rect 549 24 552 25
rect 566 27 576 31
rect 531 23 554 24
rect 560 23 576 27
rect 531 0 576 23
rect 579 42 589 45
rect 579 36 585 42
rect 597 40 599 43
rect 601 40 609 43
rect 611 40 612 43
rect 579 34 588 36
rect 735 50 736 53
rect 738 50 746 53
rect 748 50 750 53
rect 762 51 768 57
rect 758 48 768 51
rect 771 70 816 93
rect 771 66 787 70
rect 793 69 816 70
rect 771 62 781 66
rect 795 68 798 69
rect 795 65 798 66
rect 771 59 782 62
rect 784 59 785 62
rect 771 57 780 59
rect 771 51 777 57
rect 803 61 816 69
rect 819 70 864 93
rect 819 69 842 70
rect 819 61 832 69
rect 837 68 840 69
rect 837 65 840 66
rect 848 66 864 70
rect 854 62 864 66
rect 803 59 814 61
rect 821 60 832 61
rect 824 59 832 60
rect 850 59 851 62
rect 853 59 864 62
rect 855 57 864 59
rect 771 48 781 51
rect 789 50 791 53
rect 793 50 801 53
rect 803 50 804 53
rect 639 40 640 43
rect 642 40 650 43
rect 652 40 654 43
rect 662 42 672 45
rect 579 31 590 34
rect 592 31 593 34
rect 611 32 622 34
rect 632 33 640 34
rect 629 32 640 33
rect 579 27 589 31
rect 579 23 595 27
rect 603 27 606 28
rect 603 24 606 25
rect 611 24 624 32
rect 601 23 624 24
rect 579 0 624 23
rect 627 24 640 32
rect 666 36 672 42
rect 663 34 672 36
rect 658 31 659 34
rect 661 31 672 34
rect 645 27 648 28
rect 645 24 648 25
rect 662 27 672 31
rect 627 23 650 24
rect 656 23 672 27
rect 627 0 672 23
rect 675 42 685 45
rect 675 36 681 42
rect 693 40 695 43
rect 697 40 705 43
rect 707 40 708 43
rect 675 34 684 36
rect 831 50 832 53
rect 834 50 842 53
rect 844 50 846 53
rect 858 51 864 57
rect 854 48 864 51
rect 867 70 912 93
rect 867 66 883 70
rect 889 69 912 70
rect 867 62 877 66
rect 891 68 894 69
rect 891 65 894 66
rect 867 59 878 62
rect 880 59 881 62
rect 867 57 876 59
rect 867 51 873 57
rect 899 61 912 69
rect 915 70 960 93
rect 915 69 938 70
rect 915 61 928 69
rect 933 68 936 69
rect 933 65 936 66
rect 944 66 960 70
rect 950 62 960 66
rect 899 59 910 61
rect 917 60 928 61
rect 920 59 928 60
rect 946 59 947 62
rect 949 59 960 62
rect 951 57 960 59
rect 867 48 877 51
rect 885 50 887 53
rect 889 50 897 53
rect 899 50 900 53
rect 735 40 736 43
rect 738 40 746 43
rect 748 40 750 43
rect 758 42 768 45
rect 675 31 686 34
rect 688 31 689 34
rect 707 32 718 34
rect 728 33 736 34
rect 725 32 736 33
rect 675 27 685 31
rect 675 23 691 27
rect 699 27 702 28
rect 699 24 702 25
rect 707 24 720 32
rect 697 23 720 24
rect 675 0 720 23
rect 723 24 736 32
rect 762 36 768 42
rect 759 34 768 36
rect 754 31 755 34
rect 757 31 768 34
rect 741 27 744 28
rect 741 24 744 25
rect 758 27 768 31
rect 723 23 746 24
rect 752 23 768 27
rect 723 0 768 23
rect 771 42 781 45
rect 771 36 777 42
rect 789 40 791 43
rect 793 40 801 43
rect 803 40 804 43
rect 771 34 780 36
rect 927 50 928 53
rect 930 50 938 53
rect 940 50 942 53
rect 954 51 960 57
rect 950 48 960 51
rect 831 40 832 43
rect 834 40 842 43
rect 844 40 846 43
rect 854 42 864 45
rect 771 31 782 34
rect 784 31 785 34
rect 803 32 814 34
rect 824 33 832 34
rect 821 32 832 33
rect 771 27 781 31
rect 771 23 787 27
rect 795 27 798 28
rect 795 24 798 25
rect 803 24 816 32
rect 793 23 816 24
rect 771 0 816 23
rect 819 24 832 32
rect 858 36 864 42
rect 855 34 864 36
rect 850 31 851 34
rect 853 31 864 34
rect 837 27 840 28
rect 837 24 840 25
rect 854 27 864 31
rect 819 23 842 24
rect 848 23 864 27
rect 819 0 864 23
rect 867 42 877 45
rect 867 36 873 42
rect 885 40 887 43
rect 889 40 897 43
rect 899 40 900 43
rect 867 34 876 36
rect 927 40 928 43
rect 930 40 938 43
rect 940 40 942 43
rect 950 42 960 45
rect 867 31 878 34
rect 880 31 881 34
rect 899 32 910 34
rect 920 33 928 34
rect 917 32 928 33
rect 867 27 877 31
rect 867 23 883 27
rect 891 27 894 28
rect 891 24 894 25
rect 899 24 912 32
rect 889 23 912 24
rect 867 0 912 23
rect 915 24 928 32
rect 954 36 960 42
rect 951 34 960 36
rect 946 31 947 34
rect 949 31 960 34
rect 933 27 936 28
rect 933 24 936 25
rect 950 27 960 31
rect 915 23 938 24
rect 944 23 960 27
rect 915 0 960 23
rect 36 -16 37 -13
rect 39 -16 40 -13
rect 59 -16 60 -13
rect 62 -16 63 -13
rect 132 -16 133 -13
rect 135 -16 136 -13
rect 28 -32 29 -29
rect 31 -32 32 -29
rect 8 -40 9 -37
rect 11 -40 14 -37
rect 16 -40 17 -37
rect 36 -32 37 -29
rect 39 -32 40 -29
rect 155 -16 156 -13
rect 158 -16 159 -13
rect 228 -16 229 -13
rect 231 -16 232 -13
rect 59 -32 60 -29
rect 62 -32 63 -29
rect 67 -32 68 -29
rect 70 -32 71 -29
rect 124 -32 125 -29
rect 127 -32 128 -29
rect 82 -40 83 -37
rect 85 -40 88 -37
rect 90 -40 91 -37
rect 104 -40 105 -37
rect 107 -40 110 -37
rect 112 -40 113 -37
rect 132 -32 133 -29
rect 135 -32 136 -29
rect 251 -16 252 -13
rect 254 -16 255 -13
rect 324 -16 325 -13
rect 327 -16 328 -13
rect 155 -32 156 -29
rect 158 -32 159 -29
rect 163 -32 164 -29
rect 166 -32 167 -29
rect 220 -32 221 -29
rect 223 -32 224 -29
rect 178 -40 179 -37
rect 181 -40 184 -37
rect 186 -40 187 -37
rect 200 -40 201 -37
rect 203 -40 206 -37
rect 208 -40 209 -37
rect 228 -32 229 -29
rect 231 -32 232 -29
rect 347 -16 348 -13
rect 350 -16 351 -13
rect 420 -16 421 -13
rect 423 -16 424 -13
rect 251 -32 252 -29
rect 254 -32 255 -29
rect 259 -32 260 -29
rect 262 -32 263 -29
rect 316 -32 317 -29
rect 319 -32 320 -29
rect 274 -40 275 -37
rect 277 -40 280 -37
rect 282 -40 283 -37
rect 296 -40 297 -37
rect 299 -40 302 -37
rect 304 -40 305 -37
rect 324 -32 325 -29
rect 327 -32 328 -29
rect 443 -16 444 -13
rect 446 -16 447 -13
rect 516 -16 517 -13
rect 519 -16 520 -13
rect 347 -32 348 -29
rect 350 -32 351 -29
rect 355 -32 356 -29
rect 358 -32 359 -29
rect 412 -32 413 -29
rect 415 -32 416 -29
rect 370 -40 371 -37
rect 373 -40 376 -37
rect 378 -40 379 -37
rect 392 -40 393 -37
rect 395 -40 398 -37
rect 400 -40 401 -37
rect 420 -32 421 -29
rect 423 -32 424 -29
rect 539 -16 540 -13
rect 542 -16 543 -13
rect 612 -16 613 -13
rect 615 -16 616 -13
rect 443 -32 444 -29
rect 446 -32 447 -29
rect 451 -32 452 -29
rect 454 -32 455 -29
rect 508 -32 509 -29
rect 511 -32 512 -29
rect 466 -40 467 -37
rect 469 -40 472 -37
rect 474 -40 475 -37
rect 488 -40 489 -37
rect 491 -40 494 -37
rect 496 -40 497 -37
rect 516 -32 517 -29
rect 519 -32 520 -29
rect 635 -16 636 -13
rect 638 -16 639 -13
rect 708 -16 709 -13
rect 711 -16 712 -13
rect 539 -32 540 -29
rect 542 -32 543 -29
rect 547 -32 548 -29
rect 550 -32 551 -29
rect 604 -32 605 -29
rect 607 -32 608 -29
rect 562 -40 563 -37
rect 565 -40 568 -37
rect 570 -40 571 -37
rect 584 -40 585 -37
rect 587 -40 590 -37
rect 592 -40 593 -37
rect 612 -32 613 -29
rect 615 -32 616 -29
rect 731 -16 732 -13
rect 734 -16 735 -13
rect 804 -16 805 -13
rect 807 -16 808 -13
rect 635 -32 636 -29
rect 638 -32 639 -29
rect 643 -32 644 -29
rect 646 -32 647 -29
rect 700 -32 701 -29
rect 703 -32 704 -29
rect 658 -40 659 -37
rect 661 -40 664 -37
rect 666 -40 667 -37
rect 680 -40 681 -37
rect 683 -40 686 -37
rect 688 -40 689 -37
rect 708 -32 709 -29
rect 711 -32 712 -29
rect 827 -16 828 -13
rect 830 -16 831 -13
rect 900 -16 901 -13
rect 903 -16 904 -13
rect 731 -32 732 -29
rect 734 -32 735 -29
rect 739 -32 740 -29
rect 742 -32 743 -29
rect 796 -32 797 -29
rect 799 -32 800 -29
rect 754 -40 755 -37
rect 757 -40 760 -37
rect 762 -40 763 -37
rect 776 -40 777 -37
rect 779 -40 782 -37
rect 784 -40 785 -37
rect 804 -32 805 -29
rect 807 -32 808 -29
rect 923 -16 924 -13
rect 926 -16 927 -13
rect 827 -32 828 -29
rect 830 -32 831 -29
rect 835 -32 836 -29
rect 838 -32 839 -29
rect 892 -32 893 -29
rect 895 -32 896 -29
rect 850 -40 851 -37
rect 853 -40 856 -37
rect 858 -40 859 -37
rect 872 -40 873 -37
rect 875 -40 878 -37
rect 880 -40 881 -37
rect 900 -32 901 -29
rect 903 -32 904 -29
rect 923 -32 924 -29
rect 926 -32 927 -29
rect 931 -32 932 -29
rect 934 -32 935 -29
rect 946 -40 947 -37
rect 949 -40 952 -37
rect 954 -40 955 -37
<< pdiffusion >>
rect 11 -16 12 -13
rect 14 -16 15 -13
rect 84 -16 85 -13
rect 87 -16 88 -13
rect 107 -16 108 -13
rect 110 -16 111 -13
rect 180 -16 181 -13
rect 183 -16 184 -13
rect 203 -16 204 -13
rect 206 -16 207 -13
rect 276 -16 277 -13
rect 279 -16 280 -13
rect 299 -16 300 -13
rect 302 -16 303 -13
rect 372 -16 373 -13
rect 375 -16 376 -13
rect 395 -16 396 -13
rect 398 -16 399 -13
rect 468 -16 469 -13
rect 471 -16 472 -13
rect 491 -16 492 -13
rect 494 -16 495 -13
rect 564 -16 565 -13
rect 567 -16 568 -13
rect 587 -16 588 -13
rect 590 -16 591 -13
rect 660 -16 661 -13
rect 663 -16 664 -13
rect 683 -16 684 -13
rect 686 -16 687 -13
rect 756 -16 757 -13
rect 759 -16 760 -13
rect 779 -16 780 -13
rect 782 -16 783 -13
rect 852 -16 853 -13
rect 855 -16 856 -13
rect 875 -16 876 -13
rect 878 -16 879 -13
rect 948 -16 949 -13
rect 951 -16 952 -13
<< ndcontact >>
rect 17 58 21 62
rect 27 61 31 65
rect 68 61 72 65
rect 78 58 82 62
rect 17 49 21 53
rect 36 49 40 53
rect 59 49 63 53
rect 78 49 82 53
rect 113 58 117 62
rect 123 61 127 65
rect 164 61 168 65
rect 174 58 178 62
rect 113 49 117 53
rect 132 49 136 53
rect 17 40 21 44
rect 36 40 40 44
rect 155 49 159 53
rect 174 49 178 53
rect 209 58 213 62
rect 219 61 223 65
rect 260 61 264 65
rect 270 58 274 62
rect 209 49 213 53
rect 228 49 232 53
rect 59 40 63 44
rect 78 40 82 44
rect 17 31 21 35
rect 27 28 31 32
rect 68 28 72 32
rect 78 31 82 35
rect 113 40 117 44
rect 132 40 136 44
rect 251 49 255 53
rect 270 49 274 53
rect 305 58 309 62
rect 315 61 319 65
rect 356 61 360 65
rect 366 58 370 62
rect 305 49 309 53
rect 324 49 328 53
rect 155 40 159 44
rect 174 40 178 44
rect 113 31 117 35
rect 123 28 127 32
rect 164 28 168 32
rect 174 31 178 35
rect 209 40 213 44
rect 228 40 232 44
rect 347 49 351 53
rect 366 49 370 53
rect 401 58 405 62
rect 411 61 415 65
rect 452 61 456 65
rect 462 58 466 62
rect 401 49 405 53
rect 420 49 424 53
rect 251 40 255 44
rect 270 40 274 44
rect 209 31 213 35
rect 219 28 223 32
rect 260 28 264 32
rect 270 31 274 35
rect 305 40 309 44
rect 324 40 328 44
rect 443 49 447 53
rect 462 49 466 53
rect 497 58 501 62
rect 507 61 511 65
rect 548 61 552 65
rect 558 58 562 62
rect 497 49 501 53
rect 516 49 520 53
rect 347 40 351 44
rect 366 40 370 44
rect 305 31 309 35
rect 315 28 319 32
rect 356 28 360 32
rect 366 31 370 35
rect 401 40 405 44
rect 420 40 424 44
rect 539 49 543 53
rect 558 49 562 53
rect 593 58 597 62
rect 603 61 607 65
rect 644 61 648 65
rect 654 58 658 62
rect 593 49 597 53
rect 612 49 616 53
rect 443 40 447 44
rect 462 40 466 44
rect 401 31 405 35
rect 411 28 415 32
rect 452 28 456 32
rect 462 31 466 35
rect 497 40 501 44
rect 516 40 520 44
rect 635 49 639 53
rect 654 49 658 53
rect 689 58 693 62
rect 699 61 703 65
rect 740 61 744 65
rect 750 58 754 62
rect 689 49 693 53
rect 708 49 712 53
rect 539 40 543 44
rect 558 40 562 44
rect 497 31 501 35
rect 507 28 511 32
rect 548 28 552 32
rect 558 31 562 35
rect 593 40 597 44
rect 612 40 616 44
rect 731 49 735 53
rect 750 49 754 53
rect 785 58 789 62
rect 795 61 799 65
rect 836 61 840 65
rect 846 58 850 62
rect 785 49 789 53
rect 804 49 808 53
rect 635 40 639 44
rect 654 40 658 44
rect 593 31 597 35
rect 603 28 607 32
rect 644 28 648 32
rect 654 31 658 35
rect 689 40 693 44
rect 708 40 712 44
rect 827 49 831 53
rect 846 49 850 53
rect 881 58 885 62
rect 891 61 895 65
rect 932 61 936 65
rect 942 58 946 62
rect 881 49 885 53
rect 900 49 904 53
rect 731 40 735 44
rect 750 40 754 44
rect 689 31 693 35
rect 699 28 703 32
rect 740 28 744 32
rect 750 31 754 35
rect 785 40 789 44
rect 804 40 808 44
rect 923 49 927 53
rect 942 49 946 53
rect 827 40 831 44
rect 846 40 850 44
rect 785 31 789 35
rect 795 28 799 32
rect 836 28 840 32
rect 846 31 850 35
rect 881 40 885 44
rect 900 40 904 44
rect 923 40 927 44
rect 942 40 946 44
rect 881 31 885 35
rect 891 28 895 32
rect 932 28 936 32
rect 942 31 946 35
rect 32 -17 36 -13
rect 40 -17 44 -13
rect 55 -17 59 -13
rect 63 -17 67 -13
rect 128 -17 132 -13
rect 24 -33 28 -29
rect 4 -41 8 -37
rect 17 -41 21 -37
rect 32 -33 36 -29
rect 40 -33 44 -29
rect 136 -17 140 -13
rect 151 -17 155 -13
rect 159 -17 163 -13
rect 224 -17 228 -13
rect 55 -33 59 -29
rect 63 -33 67 -29
rect 71 -33 75 -29
rect 120 -33 124 -29
rect 78 -41 82 -37
rect 91 -41 95 -37
rect 100 -41 104 -37
rect 113 -41 117 -37
rect 128 -33 132 -29
rect 136 -33 140 -29
rect 232 -17 236 -13
rect 247 -17 251 -13
rect 255 -17 259 -13
rect 320 -17 324 -13
rect 151 -33 155 -29
rect 159 -33 163 -29
rect 167 -33 171 -29
rect 216 -33 220 -29
rect 174 -41 178 -37
rect 187 -41 191 -37
rect 196 -41 200 -37
rect 209 -41 213 -37
rect 224 -33 228 -29
rect 232 -33 236 -29
rect 328 -17 332 -13
rect 343 -17 347 -13
rect 351 -17 355 -13
rect 416 -17 420 -13
rect 247 -33 251 -29
rect 255 -33 259 -29
rect 263 -33 267 -29
rect 312 -33 316 -29
rect 270 -41 274 -37
rect 283 -41 287 -37
rect 292 -41 296 -37
rect 305 -41 309 -37
rect 320 -33 324 -29
rect 328 -33 332 -29
rect 424 -17 428 -13
rect 439 -17 443 -13
rect 447 -17 451 -13
rect 512 -17 516 -13
rect 343 -33 347 -29
rect 351 -33 355 -29
rect 359 -33 363 -29
rect 408 -33 412 -29
rect 366 -41 370 -37
rect 379 -41 383 -37
rect 388 -41 392 -37
rect 401 -41 405 -37
rect 416 -33 420 -29
rect 424 -33 428 -29
rect 520 -17 524 -13
rect 535 -17 539 -13
rect 543 -17 547 -13
rect 608 -17 612 -13
rect 439 -33 443 -29
rect 447 -33 451 -29
rect 455 -33 459 -29
rect 504 -33 508 -29
rect 462 -41 466 -37
rect 475 -41 479 -37
rect 484 -41 488 -37
rect 497 -41 501 -37
rect 512 -33 516 -29
rect 520 -33 524 -29
rect 616 -17 620 -13
rect 631 -17 635 -13
rect 639 -17 643 -13
rect 704 -17 708 -13
rect 535 -33 539 -29
rect 543 -33 547 -29
rect 551 -33 555 -29
rect 600 -33 604 -29
rect 558 -41 562 -37
rect 571 -41 575 -37
rect 580 -41 584 -37
rect 593 -41 597 -37
rect 608 -33 612 -29
rect 616 -33 620 -29
rect 712 -17 716 -13
rect 727 -17 731 -13
rect 735 -17 739 -13
rect 800 -17 804 -13
rect 631 -33 635 -29
rect 639 -33 643 -29
rect 647 -33 651 -29
rect 696 -33 700 -29
rect 654 -41 658 -37
rect 667 -41 671 -37
rect 676 -41 680 -37
rect 689 -41 693 -37
rect 704 -33 708 -29
rect 712 -33 716 -29
rect 808 -17 812 -13
rect 823 -17 827 -13
rect 831 -17 835 -13
rect 896 -17 900 -13
rect 727 -33 731 -29
rect 735 -33 739 -29
rect 743 -33 747 -29
rect 792 -33 796 -29
rect 750 -41 754 -37
rect 763 -41 767 -37
rect 772 -41 776 -37
rect 785 -41 789 -37
rect 800 -33 804 -29
rect 808 -33 812 -29
rect 904 -17 908 -13
rect 919 -17 923 -13
rect 927 -17 931 -13
rect 823 -33 827 -29
rect 831 -33 835 -29
rect 839 -33 843 -29
rect 888 -33 892 -29
rect 846 -41 850 -37
rect 859 -41 863 -37
rect 868 -41 872 -37
rect 881 -41 885 -37
rect 896 -33 900 -29
rect 904 -33 908 -29
rect 919 -33 923 -29
rect 927 -33 931 -29
rect 935 -33 939 -29
rect 942 -41 946 -37
rect 955 -41 959 -37
<< pdcontact >>
rect 7 -17 11 -13
rect 15 -17 19 -13
rect 80 -17 84 -13
rect 88 -17 92 -13
rect 103 -17 107 -13
rect 111 -17 115 -13
rect 176 -17 180 -13
rect 184 -17 188 -13
rect 199 -17 203 -13
rect 207 -17 211 -13
rect 272 -17 276 -13
rect 280 -17 284 -13
rect 295 -17 299 -13
rect 303 -17 307 -13
rect 368 -17 372 -13
rect 376 -17 380 -13
rect 391 -17 395 -13
rect 399 -17 403 -13
rect 464 -17 468 -13
rect 472 -17 476 -13
rect 487 -17 491 -13
rect 495 -17 499 -13
rect 560 -17 564 -13
rect 568 -17 572 -13
rect 583 -17 587 -13
rect 591 -17 595 -13
rect 656 -17 660 -13
rect 664 -17 668 -13
rect 679 -17 683 -13
rect 687 -17 691 -13
rect 752 -17 756 -13
rect 760 -17 764 -13
rect 775 -17 779 -13
rect 783 -17 787 -13
rect 848 -17 852 -13
rect 856 -17 860 -13
rect 871 -17 875 -13
rect 879 -17 883 -13
rect 944 -17 948 -13
rect 952 -17 956 -13
<< psubstratepdiff >>
rect 44 53 55 54
rect 44 47 45 53
rect 54 47 55 53
rect 140 53 151 54
rect 44 39 55 47
rect 140 47 141 53
rect 150 47 151 53
rect 236 53 247 54
rect 140 39 151 47
rect 236 47 237 53
rect 246 47 247 53
rect 332 53 343 54
rect 236 39 247 47
rect 332 47 333 53
rect 342 47 343 53
rect 428 53 439 54
rect 332 39 343 47
rect 428 47 429 53
rect 438 47 439 53
rect 524 53 535 54
rect 428 39 439 47
rect 524 47 525 53
rect 534 47 535 53
rect 620 53 631 54
rect 524 39 535 47
rect 620 47 621 53
rect 630 47 631 53
rect 716 53 727 54
rect 620 39 631 47
rect 716 47 717 53
rect 726 47 727 53
rect 812 53 823 54
rect 716 39 727 47
rect 812 47 813 53
rect 822 47 823 53
rect 908 53 919 54
rect 812 39 823 47
rect 908 47 909 53
rect 918 47 919 53
rect 908 39 919 47
<< nsubstratendiff >>
rect 0 -13 7 -12
rect 92 -13 103 -12
rect 188 -13 199 -12
rect 284 -13 295 -12
rect 380 -13 391 -12
rect 476 -13 487 -12
rect 572 -13 583 -12
rect 668 -13 679 -12
rect 764 -13 775 -12
rect 860 -13 871 -12
rect 956 -13 963 -12
rect 5 -17 7 -13
rect 0 -18 7 -17
rect 92 -17 94 -13
rect 101 -17 103 -13
rect 92 -18 103 -17
rect 188 -17 190 -13
rect 197 -17 199 -13
rect 188 -18 199 -17
rect 284 -17 286 -13
rect 293 -17 295 -13
rect 284 -18 295 -17
rect 380 -17 382 -13
rect 389 -17 391 -13
rect 380 -18 391 -17
rect 476 -17 478 -13
rect 485 -17 487 -13
rect 476 -18 487 -17
rect 572 -17 574 -13
rect 581 -17 583 -13
rect 572 -18 583 -17
rect 668 -17 670 -13
rect 677 -17 679 -13
rect 668 -18 679 -17
rect 764 -17 766 -13
rect 773 -17 775 -13
rect 764 -18 775 -17
rect 860 -17 862 -13
rect 869 -17 871 -13
rect 860 -18 871 -17
rect 956 -17 958 -13
rect 962 -17 963 -13
rect 956 -18 963 -17
<< psubstratepcontact >>
rect 45 47 54 53
rect 141 47 150 53
rect 237 47 246 53
rect 333 47 342 53
rect 429 47 438 53
rect 525 47 534 53
rect 621 47 630 53
rect 717 47 726 53
rect 813 47 822 53
rect 909 47 918 53
<< nsubstratencontact >>
rect 0 -17 5 -13
rect 94 -17 101 -13
rect 190 -17 197 -13
rect 286 -17 293 -13
rect 382 -17 389 -13
rect 478 -17 485 -13
rect 574 -17 581 -13
rect 670 -17 677 -13
rect 766 -17 773 -13
rect 862 -17 869 -13
rect 958 -17 962 -13
<< polysilicon >>
rect 24 66 27 68
rect 30 66 32 68
rect 14 62 16 64
rect 14 53 16 59
rect 67 66 69 68
rect 72 66 75 68
rect 83 62 85 64
rect 23 53 25 56
rect 33 56 47 58
rect 52 59 53 60
rect 52 58 56 59
rect 52 56 66 58
rect 33 53 35 56
rect 64 53 66 56
rect 74 53 76 56
rect 83 53 85 59
rect 23 48 25 50
rect 33 48 35 50
rect 64 48 66 50
rect 74 48 76 50
rect 120 66 123 68
rect 126 66 128 68
rect 110 62 112 64
rect 110 53 112 59
rect 163 66 165 68
rect 168 66 171 68
rect 179 62 181 64
rect 119 53 121 56
rect 129 56 143 58
rect 148 59 149 60
rect 148 58 152 59
rect 148 56 162 58
rect 129 53 131 56
rect 160 53 162 56
rect 170 53 172 56
rect 179 53 181 59
rect 119 48 121 50
rect 129 48 131 50
rect 23 43 25 45
rect 33 43 35 45
rect 14 34 16 40
rect 23 37 25 40
rect 33 37 35 40
rect 160 48 162 50
rect 170 48 172 50
rect 216 66 219 68
rect 222 66 224 68
rect 206 62 208 64
rect 206 53 208 59
rect 259 66 261 68
rect 264 66 267 68
rect 275 62 277 64
rect 215 53 217 56
rect 225 56 239 58
rect 244 59 245 60
rect 244 58 248 59
rect 244 56 258 58
rect 225 53 227 56
rect 256 53 258 56
rect 266 53 268 56
rect 275 53 277 59
rect 215 48 217 50
rect 225 48 227 50
rect 64 43 66 45
rect 74 43 76 45
rect 64 37 66 40
rect 33 35 47 37
rect 52 35 66 37
rect 74 37 76 40
rect 52 34 56 35
rect 52 33 53 34
rect 14 29 16 31
rect 24 25 27 27
rect 30 25 32 27
rect 83 34 85 40
rect 83 29 85 31
rect 67 25 69 27
rect 72 25 75 27
rect 119 43 121 45
rect 129 43 131 45
rect 110 34 112 40
rect 119 37 121 40
rect 129 37 131 40
rect 256 48 258 50
rect 266 48 268 50
rect 312 66 315 68
rect 318 66 320 68
rect 302 62 304 64
rect 302 53 304 59
rect 355 66 357 68
rect 360 66 363 68
rect 371 62 373 64
rect 311 53 313 56
rect 321 56 335 58
rect 340 59 341 60
rect 340 58 344 59
rect 340 56 354 58
rect 321 53 323 56
rect 352 53 354 56
rect 362 53 364 56
rect 371 53 373 59
rect 311 48 313 50
rect 321 48 323 50
rect 160 43 162 45
rect 170 43 172 45
rect 160 37 162 40
rect 129 35 143 37
rect 148 35 162 37
rect 170 37 172 40
rect 148 34 152 35
rect 148 33 149 34
rect 110 29 112 31
rect 120 25 123 27
rect 126 25 128 27
rect 179 34 181 40
rect 179 29 181 31
rect 163 25 165 27
rect 168 25 171 27
rect 215 43 217 45
rect 225 43 227 45
rect 206 34 208 40
rect 215 37 217 40
rect 225 37 227 40
rect 352 48 354 50
rect 362 48 364 50
rect 408 66 411 68
rect 414 66 416 68
rect 398 62 400 64
rect 398 53 400 59
rect 451 66 453 68
rect 456 66 459 68
rect 467 62 469 64
rect 407 53 409 56
rect 417 56 431 58
rect 436 59 437 60
rect 436 58 440 59
rect 436 56 450 58
rect 417 53 419 56
rect 448 53 450 56
rect 458 53 460 56
rect 467 53 469 59
rect 407 48 409 50
rect 417 48 419 50
rect 256 43 258 45
rect 266 43 268 45
rect 256 37 258 40
rect 225 35 239 37
rect 244 35 258 37
rect 266 37 268 40
rect 244 34 248 35
rect 244 33 245 34
rect 206 29 208 31
rect 216 25 219 27
rect 222 25 224 27
rect 275 34 277 40
rect 275 29 277 31
rect 259 25 261 27
rect 264 25 267 27
rect 311 43 313 45
rect 321 43 323 45
rect 302 34 304 40
rect 311 37 313 40
rect 321 37 323 40
rect 448 48 450 50
rect 458 48 460 50
rect 504 66 507 68
rect 510 66 512 68
rect 494 62 496 64
rect 494 53 496 59
rect 547 66 549 68
rect 552 66 555 68
rect 563 62 565 64
rect 503 53 505 56
rect 513 56 527 58
rect 532 59 533 60
rect 532 58 536 59
rect 532 56 546 58
rect 513 53 515 56
rect 544 53 546 56
rect 554 53 556 56
rect 563 53 565 59
rect 503 48 505 50
rect 513 48 515 50
rect 352 43 354 45
rect 362 43 364 45
rect 352 37 354 40
rect 321 35 335 37
rect 340 35 354 37
rect 362 37 364 40
rect 340 34 344 35
rect 340 33 341 34
rect 302 29 304 31
rect 312 25 315 27
rect 318 25 320 27
rect 371 34 373 40
rect 371 29 373 31
rect 355 25 357 27
rect 360 25 363 27
rect 407 43 409 45
rect 417 43 419 45
rect 398 34 400 40
rect 407 37 409 40
rect 417 37 419 40
rect 544 48 546 50
rect 554 48 556 50
rect 600 66 603 68
rect 606 66 608 68
rect 590 62 592 64
rect 590 53 592 59
rect 643 66 645 68
rect 648 66 651 68
rect 659 62 661 64
rect 599 53 601 56
rect 609 56 623 58
rect 628 59 629 60
rect 628 58 632 59
rect 628 56 642 58
rect 609 53 611 56
rect 640 53 642 56
rect 650 53 652 56
rect 659 53 661 59
rect 599 48 601 50
rect 609 48 611 50
rect 448 43 450 45
rect 458 43 460 45
rect 448 37 450 40
rect 417 35 431 37
rect 436 35 450 37
rect 458 37 460 40
rect 436 34 440 35
rect 436 33 437 34
rect 398 29 400 31
rect 408 25 411 27
rect 414 25 416 27
rect 467 34 469 40
rect 467 29 469 31
rect 451 25 453 27
rect 456 25 459 27
rect 503 43 505 45
rect 513 43 515 45
rect 494 34 496 40
rect 503 37 505 40
rect 513 37 515 40
rect 640 48 642 50
rect 650 48 652 50
rect 696 66 699 68
rect 702 66 704 68
rect 686 62 688 64
rect 686 53 688 59
rect 739 66 741 68
rect 744 66 747 68
rect 755 62 757 64
rect 695 53 697 56
rect 705 56 719 58
rect 724 59 725 60
rect 724 58 728 59
rect 724 56 738 58
rect 705 53 707 56
rect 736 53 738 56
rect 746 53 748 56
rect 755 53 757 59
rect 695 48 697 50
rect 705 48 707 50
rect 544 43 546 45
rect 554 43 556 45
rect 544 37 546 40
rect 513 35 527 37
rect 532 35 546 37
rect 554 37 556 40
rect 532 34 536 35
rect 532 33 533 34
rect 494 29 496 31
rect 504 25 507 27
rect 510 25 512 27
rect 563 34 565 40
rect 563 29 565 31
rect 547 25 549 27
rect 552 25 555 27
rect 599 43 601 45
rect 609 43 611 45
rect 590 34 592 40
rect 599 37 601 40
rect 609 37 611 40
rect 736 48 738 50
rect 746 48 748 50
rect 792 66 795 68
rect 798 66 800 68
rect 782 62 784 64
rect 782 53 784 59
rect 835 66 837 68
rect 840 66 843 68
rect 851 62 853 64
rect 791 53 793 56
rect 801 56 815 58
rect 820 59 821 60
rect 820 58 824 59
rect 820 56 834 58
rect 801 53 803 56
rect 832 53 834 56
rect 842 53 844 56
rect 851 53 853 59
rect 791 48 793 50
rect 801 48 803 50
rect 640 43 642 45
rect 650 43 652 45
rect 640 37 642 40
rect 609 35 623 37
rect 628 35 642 37
rect 650 37 652 40
rect 628 34 632 35
rect 628 33 629 34
rect 590 29 592 31
rect 600 25 603 27
rect 606 25 608 27
rect 659 34 661 40
rect 659 29 661 31
rect 643 25 645 27
rect 648 25 651 27
rect 695 43 697 45
rect 705 43 707 45
rect 686 34 688 40
rect 695 37 697 40
rect 705 37 707 40
rect 832 48 834 50
rect 842 48 844 50
rect 888 66 891 68
rect 894 66 896 68
rect 878 62 880 64
rect 878 53 880 59
rect 931 66 933 68
rect 936 66 939 68
rect 947 62 949 64
rect 887 53 889 56
rect 897 56 911 58
rect 916 59 917 60
rect 916 58 920 59
rect 916 56 930 58
rect 897 53 899 56
rect 928 53 930 56
rect 938 53 940 56
rect 947 53 949 59
rect 887 48 889 50
rect 897 48 899 50
rect 736 43 738 45
rect 746 43 748 45
rect 736 37 738 40
rect 705 35 719 37
rect 724 35 738 37
rect 746 37 748 40
rect 724 34 728 35
rect 724 33 725 34
rect 686 29 688 31
rect 696 25 699 27
rect 702 25 704 27
rect 755 34 757 40
rect 755 29 757 31
rect 739 25 741 27
rect 744 25 747 27
rect 791 43 793 45
rect 801 43 803 45
rect 782 34 784 40
rect 791 37 793 40
rect 801 37 803 40
rect 928 48 930 50
rect 938 48 940 50
rect 832 43 834 45
rect 842 43 844 45
rect 832 37 834 40
rect 801 35 815 37
rect 820 35 834 37
rect 842 37 844 40
rect 820 34 824 35
rect 820 33 821 34
rect 782 29 784 31
rect 792 25 795 27
rect 798 25 800 27
rect 851 34 853 40
rect 851 29 853 31
rect 835 25 837 27
rect 840 25 843 27
rect 887 43 889 45
rect 897 43 899 45
rect 878 34 880 40
rect 887 37 889 40
rect 897 37 899 40
rect 928 43 930 45
rect 938 43 940 45
rect 928 37 930 40
rect 897 35 911 37
rect 916 35 930 37
rect 938 37 940 40
rect 916 34 920 35
rect 916 33 917 34
rect 878 29 880 31
rect 888 25 891 27
rect 894 25 896 27
rect 947 34 949 40
rect 947 29 949 31
rect 931 25 933 27
rect 936 25 939 27
rect 12 -13 14 -10
rect 37 -13 39 -11
rect 60 -13 62 -11
rect 85 -13 87 -10
rect 108 -13 110 -10
rect 133 -13 135 -11
rect 156 -13 158 -11
rect 181 -13 183 -10
rect 204 -13 206 -10
rect 229 -13 231 -11
rect 252 -13 254 -11
rect 277 -13 279 -10
rect 300 -13 302 -10
rect 325 -13 327 -11
rect 348 -13 350 -11
rect 373 -13 375 -10
rect 396 -13 398 -10
rect 421 -13 423 -11
rect 444 -13 446 -11
rect 469 -13 471 -10
rect 492 -13 494 -10
rect 517 -13 519 -11
rect 540 -13 542 -11
rect 565 -13 567 -10
rect 588 -13 590 -10
rect 613 -13 615 -11
rect 636 -13 638 -11
rect 661 -13 663 -10
rect 684 -13 686 -10
rect 709 -13 711 -11
rect 732 -13 734 -11
rect 757 -13 759 -10
rect 780 -13 782 -10
rect 805 -13 807 -11
rect 828 -13 830 -11
rect 853 -13 855 -10
rect 876 -13 878 -10
rect 901 -13 903 -11
rect 924 -13 926 -11
rect 949 -13 951 -10
rect 12 -18 14 -16
rect 37 -21 39 -16
rect 60 -21 62 -16
rect 85 -18 87 -16
rect 108 -18 110 -16
rect 37 -23 48 -21
rect 10 -27 11 -25
rect 9 -37 11 -27
rect 14 -27 15 -25
rect 14 -37 16 -27
rect 29 -28 39 -26
rect 29 -29 31 -28
rect 37 -29 39 -28
rect 9 -42 11 -40
rect 14 -42 16 -40
rect 29 -44 31 -32
rect 37 -34 39 -32
rect 46 -48 48 -23
rect 41 -49 48 -48
rect 45 -50 48 -49
rect 51 -23 62 -21
rect 133 -21 135 -16
rect 156 -21 158 -16
rect 181 -18 183 -16
rect 204 -18 206 -16
rect 133 -23 144 -21
rect 51 -48 53 -23
rect 60 -28 70 -26
rect 84 -27 85 -25
rect 60 -29 62 -28
rect 68 -29 70 -28
rect 60 -34 62 -32
rect 68 -44 70 -32
rect 83 -37 85 -27
rect 88 -27 89 -25
rect 106 -27 107 -25
rect 88 -37 90 -27
rect 105 -37 107 -27
rect 110 -27 111 -25
rect 110 -37 112 -27
rect 125 -28 135 -26
rect 125 -29 127 -28
rect 133 -29 135 -28
rect 83 -42 85 -40
rect 88 -42 90 -40
rect 105 -42 107 -40
rect 110 -42 112 -40
rect 125 -44 127 -32
rect 133 -34 135 -32
rect 142 -48 144 -23
rect 51 -49 58 -48
rect 51 -50 54 -49
rect 137 -49 144 -48
rect 141 -50 144 -49
rect 147 -23 158 -21
rect 229 -21 231 -16
rect 252 -21 254 -16
rect 277 -18 279 -16
rect 300 -18 302 -16
rect 229 -23 240 -21
rect 147 -48 149 -23
rect 156 -28 166 -26
rect 180 -27 181 -25
rect 156 -29 158 -28
rect 164 -29 166 -28
rect 156 -34 158 -32
rect 164 -44 166 -32
rect 179 -37 181 -27
rect 184 -27 185 -25
rect 202 -27 203 -25
rect 184 -37 186 -27
rect 201 -37 203 -27
rect 206 -27 207 -25
rect 206 -37 208 -27
rect 221 -28 231 -26
rect 221 -29 223 -28
rect 229 -29 231 -28
rect 179 -42 181 -40
rect 184 -42 186 -40
rect 201 -42 203 -40
rect 206 -42 208 -40
rect 221 -44 223 -32
rect 229 -34 231 -32
rect 238 -48 240 -23
rect 147 -49 154 -48
rect 147 -50 150 -49
rect 233 -49 240 -48
rect 237 -50 240 -49
rect 243 -23 254 -21
rect 325 -21 327 -16
rect 348 -21 350 -16
rect 373 -18 375 -16
rect 396 -18 398 -16
rect 325 -23 336 -21
rect 243 -48 245 -23
rect 252 -28 262 -26
rect 276 -27 277 -25
rect 252 -29 254 -28
rect 260 -29 262 -28
rect 252 -34 254 -32
rect 260 -44 262 -32
rect 275 -37 277 -27
rect 280 -27 281 -25
rect 298 -27 299 -25
rect 280 -37 282 -27
rect 297 -37 299 -27
rect 302 -27 303 -25
rect 302 -37 304 -27
rect 317 -28 327 -26
rect 317 -29 319 -28
rect 325 -29 327 -28
rect 275 -42 277 -40
rect 280 -42 282 -40
rect 297 -42 299 -40
rect 302 -42 304 -40
rect 317 -44 319 -32
rect 325 -34 327 -32
rect 334 -48 336 -23
rect 243 -49 250 -48
rect 243 -50 246 -49
rect 329 -49 336 -48
rect 333 -50 336 -49
rect 339 -23 350 -21
rect 421 -21 423 -16
rect 444 -21 446 -16
rect 469 -18 471 -16
rect 492 -18 494 -16
rect 421 -23 432 -21
rect 339 -48 341 -23
rect 348 -28 358 -26
rect 372 -27 373 -25
rect 348 -29 350 -28
rect 356 -29 358 -28
rect 348 -34 350 -32
rect 356 -44 358 -32
rect 371 -37 373 -27
rect 376 -27 377 -25
rect 394 -27 395 -25
rect 376 -37 378 -27
rect 393 -37 395 -27
rect 398 -27 399 -25
rect 398 -37 400 -27
rect 413 -28 423 -26
rect 413 -29 415 -28
rect 421 -29 423 -28
rect 371 -42 373 -40
rect 376 -42 378 -40
rect 393 -42 395 -40
rect 398 -42 400 -40
rect 413 -44 415 -32
rect 421 -34 423 -32
rect 430 -48 432 -23
rect 339 -49 346 -48
rect 339 -50 342 -49
rect 425 -49 432 -48
rect 429 -50 432 -49
rect 435 -23 446 -21
rect 517 -21 519 -16
rect 540 -21 542 -16
rect 565 -18 567 -16
rect 588 -18 590 -16
rect 517 -23 528 -21
rect 435 -48 437 -23
rect 444 -28 454 -26
rect 468 -27 469 -25
rect 444 -29 446 -28
rect 452 -29 454 -28
rect 444 -34 446 -32
rect 452 -44 454 -32
rect 467 -37 469 -27
rect 472 -27 473 -25
rect 490 -27 491 -25
rect 472 -37 474 -27
rect 489 -37 491 -27
rect 494 -27 495 -25
rect 494 -37 496 -27
rect 509 -28 519 -26
rect 509 -29 511 -28
rect 517 -29 519 -28
rect 467 -42 469 -40
rect 472 -42 474 -40
rect 489 -42 491 -40
rect 494 -42 496 -40
rect 509 -44 511 -32
rect 517 -34 519 -32
rect 526 -48 528 -23
rect 435 -49 442 -48
rect 435 -50 438 -49
rect 521 -49 528 -48
rect 525 -50 528 -49
rect 531 -23 542 -21
rect 613 -21 615 -16
rect 636 -21 638 -16
rect 661 -18 663 -16
rect 684 -18 686 -16
rect 613 -23 624 -21
rect 531 -48 533 -23
rect 540 -28 550 -26
rect 564 -27 565 -25
rect 540 -29 542 -28
rect 548 -29 550 -28
rect 540 -34 542 -32
rect 548 -44 550 -32
rect 563 -37 565 -27
rect 568 -27 569 -25
rect 586 -27 587 -25
rect 568 -37 570 -27
rect 585 -37 587 -27
rect 590 -27 591 -25
rect 590 -37 592 -27
rect 605 -28 615 -26
rect 605 -29 607 -28
rect 613 -29 615 -28
rect 563 -42 565 -40
rect 568 -42 570 -40
rect 585 -42 587 -40
rect 590 -42 592 -40
rect 605 -44 607 -32
rect 613 -34 615 -32
rect 622 -48 624 -23
rect 531 -49 538 -48
rect 531 -50 534 -49
rect 617 -49 624 -48
rect 621 -50 624 -49
rect 627 -23 638 -21
rect 709 -21 711 -16
rect 732 -21 734 -16
rect 757 -18 759 -16
rect 780 -18 782 -16
rect 709 -23 720 -21
rect 627 -48 629 -23
rect 636 -28 646 -26
rect 660 -27 661 -25
rect 636 -29 638 -28
rect 644 -29 646 -28
rect 636 -34 638 -32
rect 644 -44 646 -32
rect 659 -37 661 -27
rect 664 -27 665 -25
rect 682 -27 683 -25
rect 664 -37 666 -27
rect 681 -37 683 -27
rect 686 -27 687 -25
rect 686 -37 688 -27
rect 701 -28 711 -26
rect 701 -29 703 -28
rect 709 -29 711 -28
rect 659 -42 661 -40
rect 664 -42 666 -40
rect 681 -42 683 -40
rect 686 -42 688 -40
rect 701 -44 703 -32
rect 709 -34 711 -32
rect 718 -48 720 -23
rect 627 -49 634 -48
rect 627 -50 630 -49
rect 713 -49 720 -48
rect 717 -50 720 -49
rect 723 -23 734 -21
rect 805 -21 807 -16
rect 828 -21 830 -16
rect 853 -18 855 -16
rect 876 -18 878 -16
rect 805 -23 816 -21
rect 723 -48 725 -23
rect 732 -28 742 -26
rect 756 -27 757 -25
rect 732 -29 734 -28
rect 740 -29 742 -28
rect 732 -34 734 -32
rect 740 -44 742 -32
rect 755 -37 757 -27
rect 760 -27 761 -25
rect 778 -27 779 -25
rect 760 -37 762 -27
rect 777 -37 779 -27
rect 782 -27 783 -25
rect 782 -37 784 -27
rect 797 -28 807 -26
rect 797 -29 799 -28
rect 805 -29 807 -28
rect 755 -42 757 -40
rect 760 -42 762 -40
rect 777 -42 779 -40
rect 782 -42 784 -40
rect 797 -44 799 -32
rect 805 -34 807 -32
rect 814 -48 816 -23
rect 723 -49 730 -48
rect 723 -50 726 -49
rect 809 -49 816 -48
rect 813 -50 816 -49
rect 819 -23 830 -21
rect 901 -21 903 -16
rect 924 -21 926 -16
rect 949 -18 951 -16
rect 901 -23 912 -21
rect 819 -48 821 -23
rect 828 -28 838 -26
rect 852 -27 853 -25
rect 828 -29 830 -28
rect 836 -29 838 -28
rect 828 -34 830 -32
rect 836 -44 838 -32
rect 851 -37 853 -27
rect 856 -27 857 -25
rect 874 -27 875 -25
rect 856 -37 858 -27
rect 873 -37 875 -27
rect 878 -27 879 -25
rect 878 -37 880 -27
rect 893 -28 903 -26
rect 893 -29 895 -28
rect 901 -29 903 -28
rect 851 -42 853 -40
rect 856 -42 858 -40
rect 873 -42 875 -40
rect 878 -42 880 -40
rect 893 -44 895 -32
rect 901 -34 903 -32
rect 910 -48 912 -23
rect 819 -49 826 -48
rect 819 -50 822 -49
rect 905 -49 912 -48
rect 909 -50 912 -49
rect 915 -23 926 -21
rect 915 -48 917 -23
rect 924 -28 934 -26
rect 948 -27 949 -25
rect 924 -29 926 -28
rect 932 -29 934 -28
rect 924 -34 926 -32
rect 932 -44 934 -32
rect 947 -37 949 -27
rect 952 -27 953 -25
rect 952 -37 954 -27
rect 947 -42 949 -40
rect 952 -42 954 -40
rect 915 -49 922 -48
rect 915 -50 918 -49
<< polycontact >>
rect 20 65 24 69
rect 10 52 14 56
rect 75 65 79 69
rect 25 54 29 58
rect 47 56 52 60
rect 70 54 74 58
rect 85 52 89 56
rect 116 65 120 69
rect 106 52 110 56
rect 171 65 175 69
rect 121 54 125 58
rect 143 56 148 60
rect 166 54 170 58
rect 10 37 14 41
rect 25 35 29 39
rect 181 52 185 56
rect 212 65 216 69
rect 202 52 206 56
rect 267 65 271 69
rect 217 54 221 58
rect 239 56 244 60
rect 262 54 266 58
rect 47 33 52 37
rect 70 35 74 39
rect 20 24 24 28
rect 85 37 89 41
rect 75 24 79 28
rect 106 37 110 41
rect 121 35 125 39
rect 277 52 281 56
rect 308 65 312 69
rect 298 52 302 56
rect 363 65 367 69
rect 313 54 317 58
rect 335 56 340 60
rect 358 54 362 58
rect 143 33 148 37
rect 166 35 170 39
rect 116 24 120 28
rect 181 37 185 41
rect 171 24 175 28
rect 202 37 206 41
rect 217 35 221 39
rect 373 52 377 56
rect 404 65 408 69
rect 394 52 398 56
rect 459 65 463 69
rect 409 54 413 58
rect 431 56 436 60
rect 454 54 458 58
rect 239 33 244 37
rect 262 35 266 39
rect 212 24 216 28
rect 277 37 281 41
rect 267 24 271 28
rect 298 37 302 41
rect 313 35 317 39
rect 469 52 473 56
rect 500 65 504 69
rect 490 52 494 56
rect 555 65 559 69
rect 505 54 509 58
rect 527 56 532 60
rect 550 54 554 58
rect 335 33 340 37
rect 358 35 362 39
rect 308 24 312 28
rect 373 37 377 41
rect 363 24 367 28
rect 394 37 398 41
rect 409 35 413 39
rect 565 52 569 56
rect 596 65 600 69
rect 586 52 590 56
rect 651 65 655 69
rect 601 54 605 58
rect 623 56 628 60
rect 646 54 650 58
rect 431 33 436 37
rect 454 35 458 39
rect 404 24 408 28
rect 469 37 473 41
rect 459 24 463 28
rect 490 37 494 41
rect 505 35 509 39
rect 661 52 665 56
rect 692 65 696 69
rect 682 52 686 56
rect 747 65 751 69
rect 697 54 701 58
rect 719 56 724 60
rect 742 54 746 58
rect 527 33 532 37
rect 550 35 554 39
rect 500 24 504 28
rect 565 37 569 41
rect 555 24 559 28
rect 586 37 590 41
rect 601 35 605 39
rect 757 52 761 56
rect 788 65 792 69
rect 778 52 782 56
rect 843 65 847 69
rect 793 54 797 58
rect 815 56 820 60
rect 838 54 842 58
rect 623 33 628 37
rect 646 35 650 39
rect 596 24 600 28
rect 661 37 665 41
rect 651 24 655 28
rect 682 37 686 41
rect 697 35 701 39
rect 853 52 857 56
rect 884 65 888 69
rect 874 52 878 56
rect 939 65 943 69
rect 889 54 893 58
rect 911 56 916 60
rect 934 54 938 58
rect 719 33 724 37
rect 742 35 746 39
rect 692 24 696 28
rect 757 37 761 41
rect 747 24 751 28
rect 778 37 782 41
rect 793 35 797 39
rect 949 52 953 56
rect 815 33 820 37
rect 838 35 842 39
rect 788 24 792 28
rect 853 37 857 41
rect 843 24 847 28
rect 874 37 878 41
rect 889 35 893 39
rect 911 33 916 37
rect 934 35 938 39
rect 884 24 888 28
rect 949 37 953 41
rect 939 24 943 28
rect 12 -10 16 -6
rect 83 -10 87 -6
rect 108 -10 112 -6
rect 179 -10 183 -6
rect 204 -10 208 -6
rect 275 -10 279 -6
rect 300 -10 304 -6
rect 371 -10 375 -6
rect 396 -10 400 -6
rect 467 -10 471 -6
rect 492 -10 496 -6
rect 563 -10 567 -6
rect 588 -10 592 -6
rect 659 -10 663 -6
rect 684 -10 688 -6
rect 755 -10 759 -6
rect 780 -10 784 -6
rect 851 -10 855 -6
rect 876 -10 880 -6
rect 947 -10 951 -6
rect 6 -27 10 -23
rect 15 -27 19 -23
rect 31 -46 35 -42
rect 41 -53 45 -49
rect 80 -27 84 -23
rect 64 -46 68 -42
rect 89 -27 93 -23
rect 102 -27 106 -23
rect 111 -27 115 -23
rect 127 -46 131 -42
rect 54 -53 58 -49
rect 137 -53 141 -49
rect 176 -27 180 -23
rect 160 -46 164 -42
rect 185 -27 189 -23
rect 198 -27 202 -23
rect 207 -27 211 -23
rect 223 -46 227 -42
rect 150 -53 154 -49
rect 233 -53 237 -49
rect 272 -27 276 -23
rect 256 -46 260 -42
rect 281 -27 285 -23
rect 294 -27 298 -23
rect 303 -27 307 -23
rect 319 -46 323 -42
rect 246 -53 250 -49
rect 329 -53 333 -49
rect 368 -27 372 -23
rect 352 -46 356 -42
rect 377 -27 381 -23
rect 390 -27 394 -23
rect 399 -27 403 -23
rect 415 -46 419 -42
rect 342 -53 346 -49
rect 425 -53 429 -49
rect 464 -27 468 -23
rect 448 -46 452 -42
rect 473 -27 477 -23
rect 486 -27 490 -23
rect 495 -27 499 -23
rect 511 -46 515 -42
rect 438 -53 442 -49
rect 521 -53 525 -49
rect 560 -27 564 -23
rect 544 -46 548 -42
rect 569 -27 573 -23
rect 582 -27 586 -23
rect 591 -27 595 -23
rect 607 -46 611 -42
rect 534 -53 538 -49
rect 617 -53 621 -49
rect 656 -27 660 -23
rect 640 -46 644 -42
rect 665 -27 669 -23
rect 678 -27 682 -23
rect 687 -27 691 -23
rect 703 -46 707 -42
rect 630 -53 634 -49
rect 713 -53 717 -49
rect 752 -27 756 -23
rect 736 -46 740 -42
rect 761 -27 765 -23
rect 774 -27 778 -23
rect 783 -27 787 -23
rect 799 -46 803 -42
rect 726 -53 730 -49
rect 809 -53 813 -49
rect 848 -27 852 -23
rect 832 -46 836 -42
rect 857 -27 861 -23
rect 870 -27 874 -23
rect 879 -27 883 -23
rect 895 -46 899 -42
rect 822 -53 826 -49
rect 905 -53 909 -49
rect 944 -27 948 -23
rect 928 -46 932 -42
rect 953 -27 957 -23
rect 918 -53 922 -49
<< metal1 >>
rect 0 62 3 96
rect 37 72 41 73
rect 48 72 51 96
rect 36 69 51 72
rect 62 69 63 72
rect 0 59 17 62
rect 26 58 30 61
rect 17 53 20 58
rect 36 53 39 69
rect 60 53 63 69
rect 96 62 99 96
rect 133 72 137 73
rect 144 72 147 96
rect 132 69 147 72
rect 158 69 159 72
rect 69 58 73 61
rect 82 59 113 62
rect 79 53 82 58
rect 122 58 126 61
rect 17 44 20 49
rect 36 44 39 49
rect 49 43 54 47
rect 60 44 63 49
rect 79 44 82 49
rect 113 53 116 58
rect 132 53 135 69
rect 156 53 159 69
rect 192 62 195 96
rect 229 72 233 73
rect 240 72 243 96
rect 228 69 243 72
rect 254 69 255 72
rect 165 58 169 61
rect 178 59 209 62
rect 175 53 178 58
rect 218 58 222 61
rect 17 35 20 40
rect 0 31 17 34
rect 26 32 30 35
rect 0 0 3 31
rect 36 24 39 40
rect 60 24 63 40
rect 79 35 82 40
rect 113 44 116 49
rect 132 44 135 49
rect 145 43 150 47
rect 156 44 159 49
rect 175 44 178 49
rect 209 53 212 58
rect 228 53 231 69
rect 252 53 255 69
rect 288 62 291 96
rect 325 72 329 73
rect 336 72 339 96
rect 324 69 339 72
rect 350 69 351 72
rect 261 58 265 61
rect 274 59 305 62
rect 271 53 274 58
rect 314 58 318 61
rect 69 32 73 35
rect 113 35 116 40
rect 82 31 113 34
rect 122 32 126 35
rect 36 21 51 24
rect 37 20 41 21
rect 48 0 51 21
rect 62 21 63 24
rect 96 0 99 31
rect 132 24 135 40
rect 156 24 159 40
rect 175 35 178 40
rect 209 44 212 49
rect 228 44 231 49
rect 241 43 246 47
rect 252 44 255 49
rect 271 44 274 49
rect 305 53 308 58
rect 324 53 327 69
rect 348 53 351 69
rect 384 62 387 96
rect 421 72 425 73
rect 432 72 435 96
rect 420 69 435 72
rect 446 69 447 72
rect 357 58 361 61
rect 370 59 401 62
rect 367 53 370 58
rect 410 58 414 61
rect 165 32 169 35
rect 209 35 212 40
rect 178 31 209 34
rect 218 32 222 35
rect 132 21 147 24
rect 133 20 137 21
rect 144 0 147 21
rect 158 21 159 24
rect 192 0 195 31
rect 228 24 231 40
rect 252 24 255 40
rect 271 35 274 40
rect 305 44 308 49
rect 324 44 327 49
rect 337 43 342 47
rect 348 44 351 49
rect 367 44 370 49
rect 401 53 404 58
rect 420 53 423 69
rect 444 53 447 69
rect 480 62 483 96
rect 517 72 521 73
rect 528 72 531 96
rect 516 69 531 72
rect 542 69 543 72
rect 453 58 457 61
rect 466 59 497 62
rect 463 53 466 58
rect 506 58 510 61
rect 261 32 265 35
rect 305 35 308 40
rect 274 31 305 34
rect 314 32 318 35
rect 228 21 243 24
rect 229 20 233 21
rect 240 0 243 21
rect 254 21 255 24
rect 288 0 291 31
rect 324 24 327 40
rect 348 24 351 40
rect 367 35 370 40
rect 401 44 404 49
rect 420 44 423 49
rect 433 43 438 47
rect 444 44 447 49
rect 463 44 466 49
rect 497 53 500 58
rect 516 53 519 69
rect 540 53 543 69
rect 576 62 579 96
rect 613 72 617 73
rect 624 72 627 96
rect 612 69 627 72
rect 638 69 639 72
rect 549 58 553 61
rect 562 59 593 62
rect 559 53 562 58
rect 602 58 606 61
rect 357 32 361 35
rect 401 35 404 40
rect 370 31 401 34
rect 410 32 414 35
rect 324 21 339 24
rect 325 20 329 21
rect 336 0 339 21
rect 350 21 351 24
rect 384 0 387 31
rect 420 24 423 40
rect 444 24 447 40
rect 463 35 466 40
rect 497 44 500 49
rect 516 44 519 49
rect 529 43 534 47
rect 540 44 543 49
rect 559 44 562 49
rect 593 53 596 58
rect 612 53 615 69
rect 636 53 639 69
rect 672 62 675 96
rect 709 72 713 73
rect 720 72 723 96
rect 708 69 723 72
rect 734 69 735 72
rect 645 58 649 61
rect 658 59 689 62
rect 655 53 658 58
rect 698 58 702 61
rect 453 32 457 35
rect 497 35 500 40
rect 466 31 497 34
rect 506 32 510 35
rect 420 21 435 24
rect 421 20 425 21
rect 432 0 435 21
rect 446 21 447 24
rect 480 0 483 31
rect 516 24 519 40
rect 540 24 543 40
rect 559 35 562 40
rect 593 44 596 49
rect 612 44 615 49
rect 625 43 630 47
rect 636 44 639 49
rect 655 44 658 49
rect 689 53 692 58
rect 708 53 711 69
rect 732 53 735 69
rect 768 62 771 96
rect 805 72 809 73
rect 816 72 819 96
rect 804 69 819 72
rect 830 69 831 72
rect 741 58 745 61
rect 754 59 785 62
rect 751 53 754 58
rect 794 58 798 61
rect 549 32 553 35
rect 593 35 596 40
rect 562 31 593 34
rect 602 32 606 35
rect 516 21 531 24
rect 517 20 521 21
rect 528 0 531 21
rect 542 21 543 24
rect 576 0 579 31
rect 612 24 615 40
rect 636 24 639 40
rect 655 35 658 40
rect 689 44 692 49
rect 708 44 711 49
rect 721 43 726 47
rect 732 44 735 49
rect 751 44 754 49
rect 785 53 788 58
rect 804 53 807 69
rect 828 53 831 69
rect 864 62 867 96
rect 901 72 905 73
rect 912 72 915 96
rect 900 69 915 72
rect 926 69 927 72
rect 837 58 841 61
rect 850 59 881 62
rect 847 53 850 58
rect 890 58 894 61
rect 645 32 649 35
rect 689 35 692 40
rect 658 31 689 34
rect 698 32 702 35
rect 612 21 627 24
rect 613 20 617 21
rect 624 0 627 21
rect 638 21 639 24
rect 672 0 675 31
rect 708 24 711 40
rect 732 24 735 40
rect 751 35 754 40
rect 785 44 788 49
rect 804 44 807 49
rect 817 43 822 47
rect 828 44 831 49
rect 847 44 850 49
rect 881 53 884 58
rect 900 53 903 69
rect 924 53 927 69
rect 933 58 937 61
rect 946 59 960 62
rect 943 53 946 58
rect 741 32 745 35
rect 785 35 788 40
rect 754 31 785 34
rect 794 32 798 35
rect 708 21 723 24
rect 709 20 713 21
rect 720 0 723 21
rect 734 21 735 24
rect 768 0 771 31
rect 804 24 807 40
rect 828 24 831 40
rect 847 35 850 40
rect 881 44 884 49
rect 900 44 903 49
rect 913 43 918 47
rect 924 44 927 49
rect 943 44 946 49
rect 837 32 841 35
rect 881 35 884 40
rect 850 31 881 34
rect 890 32 894 35
rect 804 21 819 24
rect 805 20 809 21
rect 816 0 819 21
rect 830 21 831 24
rect 864 0 867 31
rect 900 24 903 40
rect 924 24 927 40
rect 943 35 946 40
rect 933 32 937 35
rect 946 31 960 34
rect 900 21 915 24
rect 901 20 905 21
rect 912 0 915 21
rect 926 21 927 24
rect 0 -3 9 0
rect 6 -13 9 -3
rect 27 -3 51 0
rect 90 -3 105 0
rect 20 -10 79 -7
rect 90 -13 93 -3
rect 102 -13 105 -3
rect 123 -3 147 0
rect 186 -3 201 0
rect 116 -10 175 -7
rect 186 -13 189 -3
rect 198 -13 201 -3
rect 219 -3 243 0
rect 282 -3 297 0
rect 212 -10 271 -7
rect 282 -13 285 -3
rect 294 -13 297 -3
rect 315 -3 339 0
rect 378 -3 393 0
rect 308 -10 367 -7
rect 378 -13 381 -3
rect 390 -13 393 -3
rect 411 -3 435 0
rect 474 -3 489 0
rect 404 -10 463 -7
rect 474 -13 477 -3
rect 486 -13 489 -3
rect 507 -3 531 0
rect 570 -3 585 0
rect 500 -10 559 -7
rect 570 -13 573 -3
rect 582 -13 585 -3
rect 603 -3 627 0
rect 666 -3 681 0
rect 596 -10 655 -7
rect 666 -13 669 -3
rect 678 -13 681 -3
rect 699 -3 723 0
rect 762 -3 777 0
rect 692 -10 751 -7
rect 762 -13 765 -3
rect 774 -13 777 -3
rect 795 -3 819 0
rect 858 -3 873 0
rect 788 -10 847 -7
rect 858 -13 861 -3
rect 870 -13 873 -3
rect 891 -3 915 0
rect 954 -3 960 0
rect 884 -10 943 -7
rect 954 -13 957 -3
rect 5 -17 7 -13
rect 19 -17 32 -13
rect 44 -16 55 -13
rect 6 -23 9 -17
rect 16 -23 19 -17
rect 19 -27 21 -23
rect 18 -37 21 -27
rect 29 -26 44 -23
rect 25 -29 28 -26
rect 41 -29 44 -26
rect 4 -44 7 -41
rect 24 -44 27 -33
rect 4 -47 27 -44
rect 24 -53 41 -50
rect 24 -56 27 -53
rect 48 -56 51 -16
rect 67 -17 80 -13
rect 92 -17 94 -13
rect 101 -17 103 -13
rect 115 -17 128 -13
rect 140 -16 151 -13
rect 55 -26 70 -23
rect 80 -23 83 -17
rect 90 -23 93 -17
rect 55 -29 58 -26
rect 71 -29 74 -26
rect 78 -27 80 -23
rect 102 -23 105 -17
rect 112 -23 115 -17
rect 115 -27 117 -23
rect 72 -44 75 -33
rect 78 -37 81 -27
rect 114 -37 117 -27
rect 125 -26 140 -23
rect 121 -29 124 -26
rect 137 -29 140 -26
rect 92 -44 95 -41
rect 72 -47 95 -44
rect 100 -44 103 -41
rect 120 -44 123 -33
rect 100 -47 123 -44
rect 58 -53 75 -50
rect 72 -56 75 -53
rect 120 -53 137 -50
rect 120 -56 123 -53
rect 144 -56 147 -16
rect 163 -17 176 -13
rect 188 -17 190 -13
rect 197 -17 199 -13
rect 211 -17 224 -13
rect 236 -16 247 -13
rect 151 -26 166 -23
rect 176 -23 179 -17
rect 186 -23 189 -17
rect 151 -29 154 -26
rect 167 -29 170 -26
rect 174 -27 176 -23
rect 198 -23 201 -17
rect 208 -23 211 -17
rect 211 -27 213 -23
rect 168 -44 171 -33
rect 174 -37 177 -27
rect 210 -37 213 -27
rect 221 -26 236 -23
rect 217 -29 220 -26
rect 233 -29 236 -26
rect 188 -44 191 -41
rect 168 -47 191 -44
rect 196 -44 199 -41
rect 216 -44 219 -33
rect 196 -47 219 -44
rect 154 -53 171 -50
rect 168 -56 171 -53
rect 216 -53 233 -50
rect 216 -56 219 -53
rect 240 -56 243 -16
rect 259 -17 272 -13
rect 284 -17 286 -13
rect 293 -17 295 -13
rect 307 -17 320 -13
rect 332 -16 343 -13
rect 247 -26 262 -23
rect 272 -23 275 -17
rect 282 -23 285 -17
rect 247 -29 250 -26
rect 263 -29 266 -26
rect 270 -27 272 -23
rect 294 -23 297 -17
rect 304 -23 307 -17
rect 307 -27 309 -23
rect 264 -44 267 -33
rect 270 -37 273 -27
rect 306 -37 309 -27
rect 317 -26 332 -23
rect 313 -29 316 -26
rect 329 -29 332 -26
rect 284 -44 287 -41
rect 264 -47 287 -44
rect 292 -44 295 -41
rect 312 -44 315 -33
rect 292 -47 315 -44
rect 250 -53 267 -50
rect 264 -56 267 -53
rect 312 -53 329 -50
rect 312 -56 315 -53
rect 336 -56 339 -16
rect 355 -17 368 -13
rect 380 -17 382 -13
rect 389 -17 391 -13
rect 403 -17 416 -13
rect 428 -16 439 -13
rect 343 -26 358 -23
rect 368 -23 371 -17
rect 378 -23 381 -17
rect 343 -29 346 -26
rect 359 -29 362 -26
rect 366 -27 368 -23
rect 390 -23 393 -17
rect 400 -23 403 -17
rect 403 -27 405 -23
rect 360 -44 363 -33
rect 366 -37 369 -27
rect 402 -37 405 -27
rect 413 -26 428 -23
rect 409 -29 412 -26
rect 425 -29 428 -26
rect 380 -44 383 -41
rect 360 -47 383 -44
rect 388 -44 391 -41
rect 408 -44 411 -33
rect 388 -47 411 -44
rect 346 -53 363 -50
rect 360 -56 363 -53
rect 408 -53 425 -50
rect 408 -56 411 -53
rect 432 -56 435 -16
rect 451 -17 464 -13
rect 476 -17 478 -13
rect 485 -17 487 -13
rect 499 -17 512 -13
rect 524 -16 535 -13
rect 439 -26 454 -23
rect 464 -23 467 -17
rect 474 -23 477 -17
rect 439 -29 442 -26
rect 455 -29 458 -26
rect 462 -27 464 -23
rect 486 -23 489 -17
rect 496 -23 499 -17
rect 499 -27 501 -23
rect 456 -44 459 -33
rect 462 -37 465 -27
rect 498 -37 501 -27
rect 509 -26 524 -23
rect 505 -29 508 -26
rect 521 -29 524 -26
rect 476 -44 479 -41
rect 456 -47 479 -44
rect 484 -44 487 -41
rect 504 -44 507 -33
rect 484 -47 507 -44
rect 442 -53 459 -50
rect 456 -56 459 -53
rect 504 -53 521 -50
rect 504 -56 507 -53
rect 528 -56 531 -16
rect 547 -17 560 -13
rect 572 -17 574 -13
rect 581 -17 583 -13
rect 595 -17 608 -13
rect 620 -16 631 -13
rect 535 -26 550 -23
rect 560 -23 563 -17
rect 570 -23 573 -17
rect 535 -29 538 -26
rect 551 -29 554 -26
rect 558 -27 560 -23
rect 582 -23 585 -17
rect 592 -23 595 -17
rect 595 -27 597 -23
rect 552 -44 555 -33
rect 558 -37 561 -27
rect 594 -37 597 -27
rect 605 -26 620 -23
rect 601 -29 604 -26
rect 617 -29 620 -26
rect 572 -44 575 -41
rect 552 -47 575 -44
rect 580 -44 583 -41
rect 600 -44 603 -33
rect 580 -47 603 -44
rect 538 -53 555 -50
rect 552 -56 555 -53
rect 600 -53 617 -50
rect 600 -56 603 -53
rect 624 -56 627 -16
rect 643 -17 656 -13
rect 668 -17 670 -13
rect 677 -17 679 -13
rect 691 -17 704 -13
rect 716 -16 727 -13
rect 631 -26 646 -23
rect 656 -23 659 -17
rect 666 -23 669 -17
rect 631 -29 634 -26
rect 647 -29 650 -26
rect 654 -27 656 -23
rect 678 -23 681 -17
rect 688 -23 691 -17
rect 691 -27 693 -23
rect 648 -44 651 -33
rect 654 -37 657 -27
rect 690 -37 693 -27
rect 701 -26 716 -23
rect 697 -29 700 -26
rect 713 -29 716 -26
rect 668 -44 671 -41
rect 648 -47 671 -44
rect 676 -44 679 -41
rect 696 -44 699 -33
rect 676 -47 699 -44
rect 634 -53 651 -50
rect 648 -56 651 -53
rect 696 -53 713 -50
rect 696 -56 699 -53
rect 720 -56 723 -16
rect 739 -17 752 -13
rect 764 -17 766 -13
rect 773 -17 775 -13
rect 787 -17 800 -13
rect 812 -16 823 -13
rect 727 -26 742 -23
rect 752 -23 755 -17
rect 762 -23 765 -17
rect 727 -29 730 -26
rect 743 -29 746 -26
rect 750 -27 752 -23
rect 774 -23 777 -17
rect 784 -23 787 -17
rect 787 -27 789 -23
rect 744 -44 747 -33
rect 750 -37 753 -27
rect 786 -37 789 -27
rect 797 -26 812 -23
rect 793 -29 796 -26
rect 809 -29 812 -26
rect 764 -44 767 -41
rect 744 -47 767 -44
rect 772 -44 775 -41
rect 792 -44 795 -33
rect 772 -47 795 -44
rect 730 -53 747 -50
rect 744 -56 747 -53
rect 792 -53 809 -50
rect 792 -56 795 -53
rect 816 -56 819 -16
rect 835 -17 848 -13
rect 860 -17 862 -13
rect 869 -17 871 -13
rect 883 -17 896 -13
rect 908 -16 919 -13
rect 823 -26 838 -23
rect 848 -23 851 -17
rect 858 -23 861 -17
rect 823 -29 826 -26
rect 839 -29 842 -26
rect 846 -27 848 -23
rect 870 -23 873 -17
rect 880 -23 883 -17
rect 883 -27 885 -23
rect 840 -44 843 -33
rect 846 -37 849 -27
rect 882 -37 885 -27
rect 893 -26 908 -23
rect 889 -29 892 -26
rect 905 -29 908 -26
rect 860 -44 863 -41
rect 840 -47 863 -44
rect 868 -44 871 -41
rect 888 -44 891 -33
rect 868 -47 891 -44
rect 826 -53 843 -50
rect 840 -56 843 -53
rect 888 -53 905 -50
rect 888 -56 891 -53
rect 912 -56 915 -16
rect 931 -17 944 -13
rect 956 -17 958 -13
rect 919 -26 934 -23
rect 944 -23 947 -17
rect 954 -23 957 -17
rect 919 -29 922 -26
rect 935 -29 938 -26
rect 942 -27 944 -23
rect 936 -44 939 -33
rect 942 -37 945 -27
rect 956 -44 959 -41
rect 936 -47 959 -44
rect 922 -53 939 -50
rect 936 -56 939 -53
<< m2contact >>
rect 58 69 62 73
rect 16 65 20 69
rect 10 48 14 52
rect 52 56 56 60
rect 79 65 83 69
rect 154 69 158 73
rect 112 65 116 69
rect 10 41 14 45
rect 45 40 49 47
rect 85 48 89 52
rect 106 48 110 52
rect 148 56 152 60
rect 175 65 179 69
rect 250 69 254 73
rect 208 65 212 69
rect 16 24 20 28
rect 52 33 56 37
rect 85 41 89 45
rect 106 41 110 45
rect 141 40 145 47
rect 181 48 185 52
rect 202 48 206 52
rect 244 56 248 60
rect 271 65 275 69
rect 346 69 350 73
rect 304 65 308 69
rect 79 24 83 28
rect 58 20 62 24
rect 112 24 116 28
rect 148 33 152 37
rect 181 41 185 45
rect 202 41 206 45
rect 237 40 241 47
rect 277 48 281 52
rect 298 48 302 52
rect 340 56 344 60
rect 367 65 371 69
rect 442 69 446 73
rect 400 65 404 69
rect 175 24 179 28
rect 154 20 158 24
rect 208 24 212 28
rect 244 33 248 37
rect 277 41 281 45
rect 298 41 302 45
rect 333 40 337 47
rect 373 48 377 52
rect 394 48 398 52
rect 436 56 440 60
rect 463 65 467 69
rect 538 69 542 73
rect 496 65 500 69
rect 271 24 275 28
rect 250 20 254 24
rect 304 24 308 28
rect 340 33 344 37
rect 373 41 377 45
rect 394 41 398 45
rect 429 40 433 47
rect 469 48 473 52
rect 490 48 494 52
rect 532 56 536 60
rect 559 65 563 69
rect 634 69 638 73
rect 592 65 596 69
rect 367 24 371 28
rect 346 20 350 24
rect 400 24 404 28
rect 436 33 440 37
rect 469 41 473 45
rect 490 41 494 45
rect 525 40 529 47
rect 565 48 569 52
rect 586 48 590 52
rect 628 56 632 60
rect 655 65 659 69
rect 730 69 734 73
rect 688 65 692 69
rect 463 24 467 28
rect 442 20 446 24
rect 496 24 500 28
rect 532 33 536 37
rect 565 41 569 45
rect 586 41 590 45
rect 621 40 625 47
rect 661 48 665 52
rect 682 48 686 52
rect 724 56 728 60
rect 751 65 755 69
rect 826 69 830 73
rect 784 65 788 69
rect 559 24 563 28
rect 538 20 542 24
rect 592 24 596 28
rect 628 33 632 37
rect 661 41 665 45
rect 682 41 686 45
rect 717 40 721 47
rect 757 48 761 52
rect 778 48 782 52
rect 820 56 824 60
rect 847 65 851 69
rect 922 69 926 73
rect 880 65 884 69
rect 655 24 659 28
rect 634 20 638 24
rect 688 24 692 28
rect 724 33 728 37
rect 757 41 761 45
rect 778 41 782 45
rect 813 40 817 47
rect 853 48 857 52
rect 874 48 878 52
rect 916 56 920 60
rect 943 65 947 69
rect 751 24 755 28
rect 730 20 734 24
rect 784 24 788 28
rect 820 33 824 37
rect 853 41 857 45
rect 874 41 878 45
rect 909 40 913 47
rect 949 48 953 52
rect 847 24 851 28
rect 826 20 830 24
rect 880 24 884 28
rect 916 33 920 37
rect 949 41 953 45
rect 943 24 947 28
rect 922 20 926 24
rect 23 -4 27 0
rect 16 -10 20 -6
rect 79 -10 83 -6
rect 119 -4 123 0
rect 112 -10 116 -6
rect 175 -10 179 -6
rect 215 -4 219 0
rect 208 -10 212 -6
rect 271 -10 275 -6
rect 311 -4 315 0
rect 304 -10 308 -6
rect 367 -10 371 -6
rect 407 -4 411 0
rect 400 -10 404 -6
rect 463 -10 467 -6
rect 503 -4 507 0
rect 496 -10 500 -6
rect 559 -10 563 -6
rect 599 -4 603 0
rect 592 -10 596 -6
rect 655 -10 659 -6
rect 695 -4 699 0
rect 688 -10 692 -6
rect 751 -10 755 -6
rect 791 -4 795 0
rect 784 -10 788 -6
rect 847 -10 851 -6
rect 887 -4 891 0
rect 880 -10 884 -6
rect 943 -10 947 -6
rect 25 -26 29 -22
rect 32 -37 36 -33
rect 35 -46 39 -42
rect 70 -26 74 -22
rect 63 -37 67 -33
rect 60 -46 64 -42
rect 121 -26 125 -22
rect 128 -37 132 -33
rect 131 -46 135 -42
rect 166 -26 170 -22
rect 159 -37 163 -33
rect 156 -46 160 -42
rect 217 -26 221 -22
rect 224 -37 228 -33
rect 227 -46 231 -42
rect 262 -26 266 -22
rect 255 -37 259 -33
rect 252 -46 256 -42
rect 313 -26 317 -22
rect 320 -37 324 -33
rect 323 -46 327 -42
rect 358 -26 362 -22
rect 351 -37 355 -33
rect 348 -46 352 -42
rect 409 -26 413 -22
rect 416 -37 420 -33
rect 419 -46 423 -42
rect 454 -26 458 -22
rect 447 -37 451 -33
rect 444 -46 448 -42
rect 505 -26 509 -22
rect 512 -37 516 -33
rect 515 -46 519 -42
rect 550 -26 554 -22
rect 543 -37 547 -33
rect 540 -46 544 -42
rect 601 -26 605 -22
rect 608 -37 612 -33
rect 611 -46 615 -42
rect 646 -26 650 -22
rect 639 -37 643 -33
rect 636 -46 640 -42
rect 697 -26 701 -22
rect 704 -37 708 -33
rect 707 -46 711 -42
rect 742 -26 746 -22
rect 735 -37 739 -33
rect 732 -46 736 -42
rect 793 -26 797 -22
rect 800 -37 804 -33
rect 803 -46 807 -42
rect 838 -26 842 -22
rect 831 -37 835 -33
rect 828 -46 832 -42
rect 889 -26 893 -22
rect 896 -37 900 -33
rect 899 -46 903 -42
rect 934 -26 938 -22
rect 927 -37 931 -33
rect 924 -46 928 -42
<< metal2 >>
rect 48 72 51 96
rect 48 69 58 72
rect 144 72 147 96
rect 144 69 154 72
rect 240 72 243 96
rect 240 69 250 72
rect 336 72 339 96
rect 336 69 346 72
rect 432 72 435 96
rect 432 69 442 72
rect 528 72 531 96
rect 528 69 538 72
rect 624 72 627 96
rect 624 69 634 72
rect 720 72 723 96
rect 720 69 730 72
rect 816 72 819 96
rect 816 69 826 72
rect 912 72 915 96
rect 912 69 922 72
rect 0 66 16 69
rect 20 66 34 69
rect 65 66 79 69
rect 31 63 68 66
rect 83 66 112 69
rect 116 66 130 69
rect 161 66 175 69
rect 127 63 164 66
rect 179 66 208 69
rect 212 66 226 69
rect 257 66 271 69
rect 223 63 260 66
rect 275 66 304 69
rect 308 66 322 69
rect 353 66 367 69
rect 319 63 356 66
rect 371 66 400 69
rect 404 66 418 69
rect 449 66 463 69
rect 415 63 452 66
rect 467 66 496 69
rect 500 66 514 69
rect 545 66 559 69
rect 511 63 548 66
rect 563 66 592 69
rect 596 66 610 69
rect 641 66 655 69
rect 607 63 644 66
rect 659 66 688 69
rect 692 66 706 69
rect 737 66 751 69
rect 703 63 740 66
rect 755 66 784 69
rect 788 66 802 69
rect 833 66 847 69
rect 799 63 836 66
rect 851 66 880 69
rect 884 66 898 69
rect 929 66 943 69
rect 895 63 932 66
rect 947 66 960 69
rect 0 59 17 62
rect 47 59 52 60
rect 14 56 52 59
rect 82 59 113 62
rect 143 59 148 60
rect 56 56 85 59
rect 110 56 148 59
rect 178 59 209 62
rect 239 59 244 60
rect 152 56 181 59
rect 206 56 244 59
rect 274 59 305 62
rect 335 59 340 60
rect 248 56 277 59
rect 302 56 340 59
rect 370 59 401 62
rect 431 59 436 60
rect 344 56 373 59
rect 398 56 436 59
rect 466 59 497 62
rect 527 59 532 60
rect 440 56 469 59
rect 494 56 532 59
rect 562 59 593 62
rect 623 59 628 60
rect 536 56 565 59
rect 590 56 628 59
rect 658 59 689 62
rect 719 59 724 60
rect 632 56 661 59
rect 686 56 724 59
rect 754 59 785 62
rect 815 59 820 60
rect 728 56 757 59
rect 782 56 820 59
rect 850 59 881 62
rect 911 59 916 60
rect 824 56 853 59
rect 878 56 916 59
rect 946 59 960 62
rect 920 56 949 59
rect 38 50 61 53
rect 38 48 41 50
rect 0 45 41 48
rect 58 48 61 50
rect 134 50 157 53
rect 134 48 137 50
rect 58 45 137 48
rect 154 48 157 50
rect 230 50 253 53
rect 230 48 233 50
rect 154 45 233 48
rect 250 48 253 50
rect 326 50 349 53
rect 326 48 329 50
rect 250 45 329 48
rect 346 48 349 50
rect 422 50 445 53
rect 422 48 425 50
rect 346 45 425 48
rect 442 48 445 50
rect 518 50 541 53
rect 518 48 521 50
rect 442 45 521 48
rect 538 48 541 50
rect 614 50 637 53
rect 614 48 617 50
rect 538 45 617 48
rect 634 48 637 50
rect 710 50 733 53
rect 710 48 713 50
rect 634 45 713 48
rect 730 48 733 50
rect 806 50 829 53
rect 806 48 809 50
rect 730 45 809 48
rect 826 48 829 50
rect 902 50 925 53
rect 902 48 905 50
rect 826 45 905 48
rect 922 48 925 50
rect 922 45 960 48
rect 14 34 52 37
rect 0 31 17 34
rect 47 33 52 34
rect 56 34 85 37
rect 110 34 148 37
rect 82 31 113 34
rect 143 33 148 34
rect 152 34 181 37
rect 206 34 244 37
rect 178 31 209 34
rect 239 33 244 34
rect 248 34 277 37
rect 302 34 340 37
rect 274 31 305 34
rect 335 33 340 34
rect 344 34 373 37
rect 398 34 436 37
rect 370 31 401 34
rect 431 33 436 34
rect 440 34 469 37
rect 494 34 532 37
rect 466 31 497 34
rect 527 33 532 34
rect 536 34 565 37
rect 590 34 628 37
rect 562 31 593 34
rect 623 33 628 34
rect 632 34 661 37
rect 686 34 724 37
rect 658 31 689 34
rect 719 33 724 34
rect 728 34 757 37
rect 782 34 820 37
rect 754 31 785 34
rect 815 33 820 34
rect 824 34 853 37
rect 878 34 916 37
rect 850 31 881 34
rect 911 33 916 34
rect 920 34 949 37
rect 946 31 960 34
rect 0 24 16 27
rect 31 27 68 30
rect 20 24 34 27
rect 65 24 79 27
rect 83 24 112 27
rect 127 27 164 30
rect 116 24 130 27
rect 161 24 175 27
rect 179 24 208 27
rect 223 27 260 30
rect 212 24 226 27
rect 257 24 271 27
rect 275 24 304 27
rect 319 27 356 30
rect 308 24 322 27
rect 353 24 367 27
rect 371 24 400 27
rect 415 27 452 30
rect 404 24 418 27
rect 449 24 463 27
rect 467 24 496 27
rect 511 27 548 30
rect 500 24 514 27
rect 545 24 559 27
rect 563 24 592 27
rect 607 27 644 30
rect 596 24 610 27
rect 641 24 655 27
rect 659 24 688 27
rect 703 27 740 30
rect 692 24 706 27
rect 737 24 751 27
rect 755 24 784 27
rect 799 27 836 30
rect 788 24 802 27
rect 833 24 847 27
rect 851 24 880 27
rect 895 27 932 30
rect 884 24 898 27
rect 929 24 943 27
rect 947 24 960 27
rect 48 21 58 24
rect 48 0 51 21
rect 144 21 154 24
rect 144 0 147 21
rect 240 21 250 24
rect 240 0 243 21
rect 336 21 346 24
rect 336 0 339 21
rect 432 21 442 24
rect 432 0 435 21
rect 528 21 538 24
rect 528 0 531 21
rect 624 21 634 24
rect 624 0 627 21
rect 720 21 730 24
rect 720 0 723 21
rect 816 21 826 24
rect 816 0 819 21
rect 912 21 922 24
rect 912 0 915 21
rect 27 -4 28 -1
rect 48 -3 74 0
rect 0 -9 16 -6
rect 12 -10 16 -9
rect 25 -22 28 -4
rect 71 -22 74 -3
rect 123 -4 124 -1
rect 144 -3 170 0
rect 83 -9 112 -6
rect 83 -10 87 -9
rect 108 -10 112 -9
rect 121 -22 124 -4
rect 167 -22 170 -3
rect 219 -4 220 -1
rect 240 -3 266 0
rect 179 -9 208 -6
rect 179 -10 183 -9
rect 204 -10 208 -9
rect 217 -22 220 -4
rect 263 -22 266 -3
rect 315 -4 316 -1
rect 336 -3 362 0
rect 275 -9 304 -6
rect 275 -10 279 -9
rect 300 -10 304 -9
rect 313 -22 316 -4
rect 359 -22 362 -3
rect 411 -4 412 -1
rect 432 -3 458 0
rect 371 -9 400 -6
rect 371 -10 375 -9
rect 396 -10 400 -9
rect 409 -22 412 -4
rect 455 -22 458 -3
rect 507 -4 508 -1
rect 528 -3 554 0
rect 467 -9 496 -6
rect 467 -10 471 -9
rect 492 -10 496 -9
rect 505 -22 508 -4
rect 551 -22 554 -3
rect 603 -4 604 -1
rect 624 -3 650 0
rect 563 -9 592 -6
rect 563 -10 567 -9
rect 588 -10 592 -9
rect 601 -22 604 -4
rect 647 -22 650 -3
rect 699 -4 700 -1
rect 720 -3 746 0
rect 659 -9 688 -6
rect 659 -10 663 -9
rect 684 -10 688 -9
rect 697 -22 700 -4
rect 743 -22 746 -3
rect 795 -4 796 -1
rect 816 -3 842 0
rect 755 -9 784 -6
rect 755 -10 759 -9
rect 780 -10 784 -9
rect 793 -22 796 -4
rect 839 -22 842 -3
rect 891 -4 892 -1
rect 912 -3 938 0
rect 851 -9 880 -6
rect 851 -10 855 -9
rect 876 -10 880 -9
rect 889 -22 892 -4
rect 935 -22 938 -3
rect 947 -9 960 -6
rect 947 -10 951 -9
rect 0 -46 35 -43
rect 39 -46 60 -43
rect 64 -46 131 -43
rect 135 -46 156 -43
rect 160 -46 227 -43
rect 231 -46 252 -43
rect 256 -46 323 -43
rect 327 -46 348 -43
rect 352 -46 419 -43
rect 423 -46 444 -43
rect 448 -46 515 -43
rect 519 -46 540 -43
rect 544 -46 611 -43
rect 615 -46 636 -43
rect 640 -46 707 -43
rect 711 -46 732 -43
rect 736 -46 803 -43
rect 807 -46 828 -43
rect 832 -46 899 -43
rect 903 -46 924 -43
rect 928 -46 960 -43
<< m3contact >>
rect 49 40 55 47
rect 145 40 151 47
rect 241 40 247 47
rect 337 40 343 47
rect 433 40 439 47
rect 529 40 535 47
rect 625 40 631 47
rect 721 40 727 47
rect 817 40 823 47
rect 913 40 919 47
rect 36 -38 40 -34
rect 59 -38 63 -34
rect 132 -38 136 -34
rect 155 -38 159 -34
rect 228 -38 232 -34
rect 251 -38 255 -34
rect 324 -38 328 -34
rect 347 -38 351 -34
rect 420 -38 424 -34
rect 443 -38 447 -34
rect 516 -38 520 -34
rect 539 -38 543 -34
rect 612 -38 616 -34
rect 635 -38 639 -34
rect 708 -38 712 -34
rect 731 -38 735 -34
rect 804 -38 808 -34
rect 827 -38 831 -34
rect 900 -38 904 -34
rect 923 -38 927 -34
<< metal3 >>
rect 13 58 35 69
rect 64 58 86 69
rect 13 49 86 58
rect 109 58 131 69
rect 160 58 182 69
rect 109 49 182 58
rect 205 58 227 69
rect 256 58 278 69
rect 205 49 278 58
rect 301 58 323 69
rect 352 58 374 69
rect 301 49 374 58
rect 397 58 419 69
rect 448 58 470 69
rect 397 49 470 58
rect 493 58 515 69
rect 544 58 566 69
rect 493 49 566 58
rect 589 58 611 69
rect 640 58 662 69
rect 589 49 662 58
rect 685 58 707 69
rect 736 58 758 69
rect 685 49 758 58
rect 781 58 803 69
rect 832 58 854 69
rect 781 49 854 58
rect 877 58 899 69
rect 928 58 950 69
rect 877 49 950 58
rect 0 47 960 49
rect 0 44 49 47
rect 13 40 49 44
rect 55 44 145 47
rect 55 40 86 44
rect 13 35 86 40
rect 13 24 35 35
rect 64 24 86 35
rect 109 40 145 44
rect 151 44 241 47
rect 151 40 182 44
rect 109 35 182 40
rect 109 24 131 35
rect 160 24 182 35
rect 205 40 241 44
rect 247 44 337 47
rect 247 40 278 44
rect 205 35 278 40
rect 205 24 227 35
rect 256 24 278 35
rect 301 40 337 44
rect 343 44 433 47
rect 343 40 374 44
rect 301 35 374 40
rect 301 24 323 35
rect 352 24 374 35
rect 397 40 433 44
rect 439 44 529 47
rect 439 40 470 44
rect 397 35 470 40
rect 397 24 419 35
rect 448 24 470 35
rect 493 40 529 44
rect 535 44 625 47
rect 535 40 566 44
rect 493 35 566 40
rect 493 24 515 35
rect 544 24 566 35
rect 589 40 625 44
rect 631 44 721 47
rect 631 40 662 44
rect 589 35 662 40
rect 589 24 611 35
rect 640 24 662 35
rect 685 40 721 44
rect 727 44 817 47
rect 727 40 758 44
rect 685 35 758 40
rect 685 24 707 35
rect 736 24 758 35
rect 781 40 817 44
rect 823 44 913 47
rect 823 40 854 44
rect 781 35 854 40
rect 781 24 803 35
rect 832 24 854 35
rect 877 40 913 44
rect 919 44 960 47
rect 919 40 950 44
rect 877 35 950 40
rect 877 24 899 35
rect 928 24 950 35
rect 35 -34 41 -33
rect 35 -38 36 -34
rect 40 -38 41 -34
rect 35 -39 41 -38
rect 58 -34 64 -33
rect 58 -38 59 -34
rect 63 -38 64 -34
rect 58 -39 64 -38
rect 131 -34 137 -33
rect 131 -38 132 -34
rect 136 -38 137 -34
rect 131 -39 137 -38
rect 154 -34 160 -33
rect 154 -38 155 -34
rect 159 -38 160 -34
rect 154 -39 160 -38
rect 227 -34 233 -33
rect 227 -38 228 -34
rect 232 -38 233 -34
rect 227 -39 233 -38
rect 250 -34 256 -33
rect 250 -38 251 -34
rect 255 -38 256 -34
rect 250 -39 256 -38
rect 323 -34 329 -33
rect 323 -38 324 -34
rect 328 -38 329 -34
rect 323 -39 329 -38
rect 346 -34 352 -33
rect 346 -38 347 -34
rect 351 -38 352 -34
rect 346 -39 352 -38
rect 419 -34 425 -33
rect 419 -38 420 -34
rect 424 -38 425 -34
rect 419 -39 425 -38
rect 442 -34 448 -33
rect 442 -38 443 -34
rect 447 -38 448 -34
rect 442 -39 448 -38
rect 515 -34 521 -33
rect 515 -38 516 -34
rect 520 -38 521 -34
rect 515 -39 521 -38
rect 538 -34 544 -33
rect 538 -38 539 -34
rect 543 -38 544 -34
rect 538 -39 544 -38
rect 611 -34 617 -33
rect 611 -38 612 -34
rect 616 -38 617 -34
rect 611 -39 617 -38
rect 634 -34 640 -33
rect 634 -38 635 -34
rect 639 -38 640 -34
rect 634 -39 640 -38
rect 707 -34 713 -33
rect 707 -38 708 -34
rect 712 -38 713 -34
rect 707 -39 713 -38
rect 730 -34 736 -33
rect 730 -38 731 -34
rect 735 -38 736 -34
rect 730 -39 736 -38
rect 803 -34 809 -33
rect 803 -38 804 -34
rect 808 -38 809 -34
rect 803 -39 809 -38
rect 826 -34 832 -33
rect 826 -38 827 -34
rect 831 -38 832 -34
rect 826 -39 832 -38
rect 899 -34 905 -33
rect 899 -38 900 -34
rect 904 -38 905 -34
rect 899 -39 905 -38
rect 922 -34 928 -33
rect 922 -38 923 -34
rect 927 -38 928 -34
rect 922 -39 928 -38
use csrldff  csrldff_0
array 0 19 48 0 0 96
timestamp 1354594767
transform 1 0 8 0 1 -152
box -13 0 35 96
<< labels >>
rlabel metal2 0 -7 0 -7 3 Vbp
rlabel metal2 96 -7 96 -7 3 Vbp
rlabel metal2 192 -7 192 -7 3 Vbp
rlabel metal2 288 -7 288 -7 3 Vbp
rlabel metal2 384 -7 384 -7 3 Vbp
rlabel metal2 480 -7 480 -7 3 Vbp
rlabel metal2 576 -7 576 -7 3 Vbp
rlabel metal2 672 -7 672 -7 3 Vbp
rlabel metal2 768 -7 768 -7 3 Vbp
rlabel metal2 864 -7 864 -7 3 Vbp
rlabel metal1 2 4 2 4 5 Vdd
rlabel metal1 98 4 98 4 5 Vdd
rlabel metal1 194 4 194 4 5 Vdd
rlabel metal1 290 4 290 4 5 Vdd
rlabel metal1 386 4 386 4 5 Vdd
rlabel metal1 482 4 482 4 5 Vdd
rlabel metal1 578 4 578 4 5 Vdd
rlabel metal1 674 4 674 4 5 Vdd
rlabel metal1 770 4 770 4 5 Vdd
rlabel metal1 866 4 866 4 5 Vdd
rlabel metal2 4 26 4 26 3 Shutter
rlabel metal2 100 26 100 26 3 Shutter
rlabel metal2 196 26 196 26 3 Shutter
rlabel metal2 292 26 292 26 3 Shutter
rlabel metal2 388 26 388 26 3 Shutter
rlabel metal2 484 26 484 26 3 Shutter
rlabel metal2 580 26 580 26 3 Shutter
rlabel metal2 676 26 676 26 3 Shutter
rlabel metal2 772 26 772 26 3 Shutter
rlabel metal2 868 26 868 26 3 Shutter
rlabel metal2 95 26 95 26 7 Shutter
rlabel metal2 191 26 191 26 7 Shutter
rlabel metal2 287 26 287 26 7 Shutter
rlabel metal2 383 26 383 26 7 Shutter
rlabel metal2 479 26 479 26 7 Shutter
rlabel metal2 575 26 575 26 7 Shutter
rlabel metal2 671 26 671 26 7 Shutter
rlabel metal2 767 26 767 26 7 Shutter
rlabel metal2 863 26 863 26 7 Shutter
rlabel metal2 959 26 959 26 7 Shutter
rlabel metal2 49 95 49 95 5 Column
rlabel metal2 145 95 145 95 5 Column
rlabel metal2 241 95 241 95 5 Column
rlabel metal2 337 95 337 95 5 Column
rlabel metal2 433 95 433 95 5 Column
rlabel metal2 529 95 529 95 5 Column
rlabel metal2 625 95 625 95 5 Column
rlabel metal2 721 95 721 95 5 Column
rlabel metal2 817 95 817 95 5 Column
rlabel metal2 913 95 913 95 5 Column
rlabel metal2 95 60 95 60 7 Row
rlabel metal2 191 60 191 60 7 Row
rlabel metal2 287 60 287 60 7 Row
rlabel metal2 383 60 383 60 7 Row
rlabel metal2 479 60 479 60 7 Row
rlabel metal2 575 60 575 60 7 Row
rlabel metal2 671 60 671 60 7 Row
rlabel metal2 767 60 767 60 7 Row
rlabel metal2 863 60 863 60 7 Row
rlabel metal2 959 60 959 60 7 Row
rlabel metal2 95 32 95 32 7 Row
rlabel metal2 191 32 191 32 7 Row
rlabel metal2 287 32 287 32 7 Row
rlabel metal2 383 32 383 32 7 Row
rlabel metal2 479 32 479 32 7 Row
rlabel metal2 575 32 575 32 7 Row
rlabel metal2 671 32 671 32 7 Row
rlabel metal2 767 32 767 32 7 Row
rlabel metal2 863 32 863 32 7 Row
rlabel metal2 959 32 959 32 7 Row
rlabel metal2 1 32 1 32 3 Row
rlabel metal2 97 32 97 32 3 Row
rlabel metal2 193 32 193 32 3 Row
rlabel metal2 289 32 289 32 3 Row
rlabel metal2 385 32 385 32 3 Row
rlabel metal2 481 32 481 32 3 Row
rlabel metal2 577 32 577 32 3 Row
rlabel metal2 673 32 673 32 3 Row
rlabel metal2 769 32 769 32 3 Row
rlabel metal2 865 32 865 32 3 Row
rlabel metal2 1 60 1 60 3 Row
rlabel metal2 97 60 97 60 3 Row
rlabel metal2 193 60 193 60 3 Row
rlabel metal2 289 60 289 60 3 Row
rlabel metal2 385 60 385 60 3 Row
rlabel metal2 481 60 481 60 3 Row
rlabel metal2 577 60 577 60 3 Row
rlabel metal2 673 60 673 60 3 Row
rlabel metal2 769 60 769 60 3 Row
rlabel metal2 865 60 865 60 3 Row
rlabel metal1 2 89 2 89 1 Vdd
rlabel metal1 98 89 98 89 1 Vdd
rlabel metal1 194 89 194 89 1 Vdd
rlabel metal1 290 89 290 89 1 Vdd
rlabel metal1 386 89 386 89 1 Vdd
rlabel metal1 482 89 482 89 1 Vdd
rlabel metal1 578 89 578 89 1 Vdd
rlabel metal1 674 89 674 89 1 Vdd
rlabel metal1 770 89 770 89 1 Vdd
rlabel metal1 866 89 866 89 1 Vdd
rlabel metal2 6 47 6 47 1 Reset
rlabel metal2 102 47 102 47 1 Reset
rlabel metal2 198 47 198 47 1 Reset
rlabel metal2 294 47 294 47 1 Reset
rlabel metal2 390 47 390 47 1 Reset
rlabel metal2 486 47 486 47 1 Reset
rlabel metal2 582 47 582 47 1 Reset
rlabel metal2 678 47 678 47 1 Reset
rlabel metal2 774 47 774 47 1 Reset
rlabel metal2 870 47 870 47 1 Reset
rlabel metal2 4 67 4 67 3 Shutter
rlabel metal2 100 67 100 67 3 Shutter
rlabel metal2 196 67 196 67 3 Shutter
rlabel metal2 292 67 292 67 3 Shutter
rlabel metal2 388 67 388 67 3 Shutter
rlabel metal2 484 67 484 67 3 Shutter
rlabel metal2 580 67 580 67 3 Shutter
rlabel metal2 676 67 676 67 3 Shutter
rlabel metal2 772 67 772 67 3 Shutter
rlabel metal2 868 67 868 67 3 Shutter
rlabel metal2 93 47 93 47 1 Reset
rlabel metal2 189 47 189 47 1 Reset
rlabel metal2 285 47 285 47 1 Reset
rlabel metal2 381 47 381 47 1 Reset
rlabel metal2 477 47 477 47 1 Reset
rlabel metal2 573 47 573 47 1 Reset
rlabel metal2 669 47 669 47 1 Reset
rlabel metal2 765 47 765 47 1 Reset
rlabel metal2 861 47 861 47 1 Reset
rlabel metal2 957 47 957 47 1 Reset
rlabel metal2 95 67 95 67 7 Shutter
rlabel metal2 191 67 191 67 7 Shutter
rlabel metal2 287 67 287 67 7 Shutter
rlabel metal2 383 67 383 67 7 Shutter
rlabel metal2 479 67 479 67 7 Shutter
rlabel metal2 575 67 575 67 7 Shutter
rlabel metal2 671 67 671 67 7 Shutter
rlabel metal2 767 67 767 67 7 Shutter
rlabel metal2 863 67 863 67 7 Shutter
rlabel metal2 959 67 959 67 7 Shutter
<< end >>
