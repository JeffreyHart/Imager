magic
tech scmos
timestamp 1354157580
<< ntransistor >>
rect -74 -39 -71 -37
rect -60 -46 -58 -43
rect -79 -56 -77 -53
rect -69 -56 -67 -53
<< ndiffusion >>
rect -89 -35 -47 -18
rect -89 -36 -69 -35
rect -89 -48 -79 -36
rect -74 -37 -71 -36
rect -74 -40 -71 -39
rect -63 -39 -47 -35
rect -57 -43 -47 -39
rect -61 -46 -60 -43
rect -58 -46 -47 -43
rect -57 -48 -47 -46
rect -80 -56 -79 -53
rect -77 -56 -69 -53
rect -67 -56 -65 -53
rect -53 -54 -47 -48
rect -57 -60 -47 -54
<< ndcontact >>
rect -75 -44 -71 -40
rect -65 -47 -61 -43
rect -84 -56 -80 -52
rect -65 -56 -61 -52
<< polysilicon >>
rect -76 -39 -74 -37
rect -71 -39 -68 -37
rect -60 -43 -58 -41
rect -79 -53 -77 -51
rect -69 -53 -67 -49
rect -60 -52 -58 -46
rect -79 -61 -77 -56
rect -69 -58 -67 -56
<< polycontact >>
rect -68 -40 -64 -36
rect -73 -51 -69 -47
rect -58 -53 -54 -49
rect -77 -62 -73 -58
<< metal1 >>
rect -92 -52 -89 -18
rect -57 -43 -54 -18
rect -74 -47 -70 -44
rect -61 -46 -54 -43
rect -64 -52 -61 -47
rect -92 -55 -84 -52
rect -92 -63 -89 -55
rect -64 -60 -61 -56
rect -64 -63 -54 -60
<< m2contact >>
rect -64 -40 -60 -36
rect -73 -63 -69 -59
rect -58 -57 -54 -53
<< metal2 >>
rect -92 -39 -64 -36
rect -60 -39 -47 -36
rect -92 -56 -58 -53
rect -54 -56 -47 -53
rect -92 -63 -73 -60
rect -69 -63 -47 -60
<< end >>
