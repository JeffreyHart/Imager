magic
tech scmos
timestamp 1354204445
use pixel  pixel_0
array 0 69 45 0 69 45
timestamp 1354157580
transform 1 0 92 0 1 63
box -92 -63 -47 -18
<< end >>
