magic
tech scmos
timestamp 1355198308
<< ntransistor >>
rect 25 -35 29 -15
rect 35 -35 39 -15
rect 45 -35 49 -15
rect 55 -35 59 -15
rect 73 -35 77 -15
rect 83 -35 87 -15
rect 93 -35 97 -15
rect 103 -35 107 -15
<< ptransistor >>
rect 5 2 9 22
rect 15 2 19 22
rect 25 2 29 22
rect 35 2 39 22
rect 45 2 49 22
rect 55 2 59 22
rect 73 2 77 22
rect 83 2 87 22
rect 93 2 97 22
rect 103 2 107 22
rect 113 2 117 22
rect 123 2 127 22
<< ndiffusion >>
rect 24 -35 25 -15
rect 29 -35 30 -15
rect 34 -35 35 -15
rect 39 -35 40 -15
rect 44 -35 45 -15
rect 49 -35 50 -15
rect 54 -35 55 -15
rect 59 -35 60 -15
rect 72 -35 73 -15
rect 77 -35 78 -15
rect 82 -35 83 -15
rect 87 -35 88 -15
rect 92 -35 93 -15
rect 97 -35 98 -15
rect 102 -35 103 -15
rect 107 -35 108 -15
<< pdiffusion >>
rect 4 2 5 22
rect 9 2 10 22
rect 14 2 15 22
rect 19 2 20 22
rect 24 2 25 22
rect 29 2 30 22
rect 34 2 35 22
rect 39 2 40 22
rect 44 2 45 22
rect 49 2 50 22
rect 54 2 55 22
rect 59 2 60 22
rect 72 2 73 22
rect 77 2 78 22
rect 82 2 83 22
rect 87 2 88 22
rect 92 2 93 22
rect 97 2 98 22
rect 102 2 103 22
rect 107 2 108 22
rect 112 2 113 22
rect 117 2 118 22
rect 122 2 123 22
rect 127 2 128 22
<< ndcontact >>
rect 20 -35 24 -15
rect 30 -35 34 -15
rect 40 -35 44 -15
rect 50 -35 54 -15
rect 60 -35 64 -15
rect 68 -35 72 -15
rect 78 -35 82 -15
rect 88 -35 92 -15
rect 98 -35 102 -15
rect 108 -35 112 -15
<< pdcontact >>
rect 0 2 4 22
rect 10 2 14 22
rect 20 2 24 22
rect 30 2 34 22
rect 40 2 44 22
rect 50 2 54 22
rect 60 2 64 22
rect 68 2 72 22
rect 78 2 82 22
rect 88 2 92 22
rect 98 2 102 22
rect 108 2 112 22
rect 118 2 122 22
rect 128 2 132 22
<< polysilicon >>
rect -1 23 19 25
rect 5 22 9 23
rect 15 22 19 23
rect 25 23 39 25
rect 25 22 29 23
rect 35 22 39 23
rect 45 23 59 25
rect 45 22 49 23
rect 55 22 59 23
rect 73 23 87 25
rect 73 22 77 23
rect 83 22 87 23
rect 93 23 107 25
rect 93 22 97 23
rect 103 22 107 23
rect 113 23 133 25
rect 113 22 117 23
rect 123 22 127 23
rect 5 0 9 2
rect 15 0 19 2
rect 25 0 29 2
rect 35 0 39 2
rect 45 0 49 2
rect 55 0 59 2
rect 25 -3 27 0
rect 0 -5 27 -3
rect 57 -4 59 0
rect 73 0 77 2
rect 83 0 87 2
rect 93 0 97 2
rect 103 0 107 2
rect 113 0 117 2
rect 123 0 127 2
rect 73 -4 75 0
rect 105 -3 107 0
rect 105 -5 132 -3
rect 25 -13 27 -9
rect 105 -13 107 -9
rect 25 -15 29 -13
rect 35 -15 39 -13
rect 45 -15 49 -13
rect 55 -15 59 -13
rect 73 -15 77 -13
rect 83 -15 87 -13
rect 93 -15 97 -13
rect 103 -15 107 -13
rect 25 -36 29 -35
rect 35 -36 39 -35
rect 45 -36 49 -35
rect 55 -36 59 -35
rect 25 -38 59 -36
rect 73 -36 77 -35
rect 83 -36 87 -35
rect 93 -36 97 -35
rect 103 -36 107 -35
rect 73 -38 107 -36
<< polycontact >>
rect 53 -4 57 0
rect 75 -4 79 0
rect 27 -13 31 -9
rect 101 -13 105 -9
<< metal1 >>
rect -1 25 14 28
rect 10 22 14 25
rect 20 25 64 28
rect 20 22 24 25
rect 40 22 44 25
rect 60 22 64 25
rect 0 -1 4 2
rect 20 -1 24 2
rect 0 -4 24 -1
rect 68 25 112 28
rect 68 22 72 25
rect 88 22 92 25
rect 108 22 112 25
rect 30 -9 34 2
rect 31 -13 34 -9
rect 30 -15 34 -13
rect 50 0 54 2
rect 78 0 82 2
rect 50 -4 53 0
rect 50 -6 57 -4
rect 79 -4 82 0
rect 50 -9 64 -6
rect 50 -15 54 -9
rect 75 -6 82 -4
rect 68 -9 82 -6
rect 78 -15 82 -9
rect 98 -9 102 2
rect 118 25 133 28
rect 118 22 122 25
rect 108 -1 112 2
rect 128 -1 132 2
rect 108 -4 132 -1
rect 98 -13 101 -9
rect 98 -15 102 -13
rect 20 -38 24 -35
rect 40 -38 44 -35
rect 60 -38 64 -35
rect -1 -41 64 -38
rect 68 -38 72 -35
rect 88 -38 92 -35
rect 108 -38 112 -35
rect 68 -41 133 -38
<< m2contact >>
rect 64 -10 68 -5
<< metal2 >>
rect 64 -5 68 28
<< labels >>
rlabel metal1 0 -40 0 -40 2 Gnd
rlabel polysilicon 0 24 0 24 4 Vb
rlabel metal1 0 27 0 27 4 Vdd
rlabel metal1 1 -4 1 -4 3 Vin
rlabel metal1 132 -40 132 -40 8 Gnd
rlabel polysilicon 132 24 132 24 6 Vb
rlabel metal1 132 27 132 27 6 Vdd
rlabel metal1 131 -4 131 -4 7 Vin
rlabel metal2 66 27 66 27 5 Vout
<< end >>
