magic
tech scmos
timestamp 1355192513
use csrldiff_vert  csrldiff_vert_1
array 0 0 113 0 31 96
timestamp 1355192033
transform 1 0 0 0 1 -2976
box -116 2967 -3 3081
use pixel_2.1  pixel_2.1_0
array 0 31 96 0 31 96
timestamp 1355189358
transform 1 0 0 0 1 0
box -3 -6 102 99
use columnamplifier  columnamplifier_0
array 0 31 96 0 0 66
timestamp 1355185946
transform 1 0 0 0 1 0
box -3 -60 102 6
use csrlend  csrlend_0
timestamp 1355186776
transform 1 0 -120 0 1 -170
box -4 7 26 87
use csrldff  csrldff_0
array 0 63 48 0 0 96
timestamp 1355188032
transform 1 0 8 0 1 -152
box -19 0 41 96
<< end >>
