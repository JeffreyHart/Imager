magic
tech scmos
timestamp 1355362639
<< nwell >>
rect 32 -24 60 -7
rect 109 -24 137 -7
<< pwell >>
rect 32 -7 137 98
rect 60 -24 109 -7
rect 32 -57 137 -24
<< ntransistor >>
rect 62 65 65 67
rect 49 58 51 61
rect 104 65 107 67
rect 88 58 91 59
rect 118 58 120 61
rect 58 49 60 52
rect 68 49 70 52
rect 99 49 101 52
rect 109 49 111 52
rect 58 39 60 42
rect 68 39 70 42
rect 99 39 101 42
rect 109 39 111 42
rect 49 30 51 33
rect 88 32 91 33
rect 62 24 65 26
rect 118 30 120 33
rect 104 24 107 26
rect 72 -17 74 -14
rect 95 -17 97 -14
rect 64 -33 66 -30
rect 44 -41 46 -38
rect 49 -41 51 -38
rect 72 -33 74 -30
rect 95 -33 97 -30
rect 103 -33 105 -30
rect 118 -41 120 -38
rect 123 -41 125 -38
<< ptransistor >>
rect 47 -17 49 -14
rect 120 -17 122 -14
<< ndiffusion >>
rect 38 69 83 92
rect 38 65 54 69
rect 60 68 83 69
rect 38 61 48 65
rect 62 67 65 68
rect 62 64 65 65
rect 38 58 49 61
rect 51 58 52 61
rect 38 56 47 58
rect 38 50 44 56
rect 70 60 83 68
rect 86 69 131 92
rect 86 68 109 69
rect 86 60 99 68
rect 104 67 107 68
rect 104 64 107 65
rect 115 65 131 69
rect 121 61 131 65
rect 70 58 81 60
rect 88 59 99 60
rect 91 58 99 59
rect 117 58 118 61
rect 120 58 131 61
rect 122 56 131 58
rect 38 47 48 50
rect 56 49 58 52
rect 60 49 68 52
rect 70 49 71 52
rect 98 49 99 52
rect 101 49 109 52
rect 111 49 113 52
rect 125 50 131 56
rect 121 47 131 50
rect 38 41 48 44
rect 38 35 44 41
rect 56 39 58 42
rect 60 39 68 42
rect 70 39 71 42
rect 38 33 47 35
rect 98 39 99 42
rect 101 39 109 42
rect 111 39 113 42
rect 121 41 131 44
rect 38 30 49 33
rect 51 30 52 33
rect 70 31 81 33
rect 91 32 99 33
rect 88 31 99 32
rect 38 26 48 30
rect 38 22 54 26
rect 62 26 65 27
rect 62 23 65 24
rect 70 23 83 31
rect 60 22 83 23
rect 38 -1 83 22
rect 86 23 99 31
rect 125 35 131 41
rect 122 33 131 35
rect 117 30 118 33
rect 120 30 131 33
rect 104 26 107 27
rect 104 23 107 24
rect 121 26 131 30
rect 86 22 109 23
rect 115 22 131 26
rect 86 -1 131 22
rect 71 -17 72 -14
rect 74 -17 75 -14
rect 94 -17 95 -14
rect 97 -17 98 -14
rect 63 -33 64 -30
rect 66 -33 67 -30
rect 43 -41 44 -38
rect 46 -41 49 -38
rect 51 -41 52 -38
rect 71 -33 72 -30
rect 74 -33 75 -30
rect 94 -33 95 -30
rect 97 -33 98 -30
rect 102 -33 103 -30
rect 105 -33 106 -30
rect 117 -41 118 -38
rect 120 -41 123 -38
rect 125 -41 126 -38
<< pdiffusion >>
rect 46 -17 47 -14
rect 49 -17 50 -14
rect 119 -17 120 -14
rect 122 -17 123 -14
<< ndcontact >>
rect 52 57 56 61
rect 62 60 66 64
rect 103 60 107 64
rect 113 57 117 61
rect 52 48 56 52
rect 71 48 75 52
rect 94 48 98 52
rect 113 48 117 52
rect 52 39 56 43
rect 71 39 75 43
rect 94 39 98 43
rect 113 39 117 43
rect 52 30 56 34
rect 62 27 66 31
rect 103 27 107 31
rect 113 30 117 34
rect 67 -18 71 -14
rect 75 -18 79 -14
rect 90 -18 94 -14
rect 98 -18 102 -14
rect 59 -34 63 -30
rect 39 -42 43 -38
rect 52 -42 56 -38
rect 67 -34 71 -30
rect 75 -34 79 -30
rect 90 -34 94 -30
rect 98 -34 102 -30
rect 106 -34 110 -30
rect 113 -42 117 -38
rect 126 -42 130 -38
<< pdcontact >>
rect 42 -18 46 -14
rect 50 -18 54 -14
rect 115 -18 119 -14
rect 123 -18 127 -14
<< psubstratepdiff >>
rect 79 52 90 53
rect 79 46 80 52
rect 89 46 90 52
rect 79 38 90 46
<< nsubstratendiff >>
rect 35 -14 42 -13
rect 127 -14 133 -13
rect 35 -18 36 -14
rect 40 -18 42 -14
rect 35 -19 42 -18
rect 127 -18 129 -14
rect 127 -19 133 -18
<< psubstratepcontact >>
rect 80 46 89 52
<< nsubstratencontact >>
rect 36 -18 40 -14
rect 129 -18 133 -14
<< polysilicon >>
rect 59 65 62 67
rect 65 65 67 67
rect 49 61 51 63
rect 49 52 51 58
rect 102 65 104 67
rect 107 65 110 67
rect 118 61 120 63
rect 58 52 60 55
rect 68 55 82 57
rect 87 58 88 59
rect 87 57 91 58
rect 87 55 101 57
rect 68 52 70 55
rect 99 52 101 55
rect 109 52 111 55
rect 118 52 120 58
rect 58 47 60 49
rect 68 47 70 49
rect 99 47 101 49
rect 109 47 111 49
rect 58 42 60 44
rect 68 42 70 44
rect 49 33 51 39
rect 58 36 60 39
rect 68 36 70 39
rect 99 42 101 44
rect 109 42 111 44
rect 99 36 101 39
rect 68 34 82 36
rect 87 34 101 36
rect 109 36 111 39
rect 87 33 91 34
rect 87 32 88 33
rect 49 28 51 30
rect 59 24 62 26
rect 65 24 67 26
rect 118 33 120 39
rect 118 28 120 30
rect 102 24 104 26
rect 107 24 110 26
rect 47 -14 49 -11
rect 72 -14 74 -12
rect 95 -14 97 -12
rect 120 -14 122 -11
rect 47 -19 49 -17
rect 72 -22 74 -17
rect 95 -22 97 -17
rect 120 -19 122 -17
rect 72 -24 83 -22
rect 45 -28 46 -26
rect 44 -38 46 -28
rect 49 -28 50 -26
rect 49 -38 51 -28
rect 64 -29 74 -27
rect 64 -30 66 -29
rect 72 -30 74 -29
rect 44 -43 46 -41
rect 49 -43 51 -41
rect 64 -45 66 -33
rect 72 -35 74 -33
rect 81 -49 83 -24
rect 76 -50 83 -49
rect 80 -51 83 -50
rect 86 -24 97 -22
rect 86 -49 88 -24
rect 95 -29 105 -27
rect 119 -28 120 -26
rect 95 -30 97 -29
rect 103 -30 105 -29
rect 95 -35 97 -33
rect 103 -45 105 -33
rect 118 -38 120 -28
rect 123 -28 124 -26
rect 123 -38 125 -28
rect 118 -43 120 -41
rect 123 -43 125 -41
rect 86 -50 93 -49
rect 86 -51 89 -50
<< polycontact >>
rect 55 64 59 68
rect 45 51 49 55
rect 110 64 114 68
rect 60 53 64 57
rect 82 55 87 59
rect 105 53 109 57
rect 120 51 124 55
rect 45 36 49 40
rect 60 34 64 38
rect 82 32 87 36
rect 105 34 109 38
rect 55 23 59 27
rect 120 36 124 40
rect 110 23 114 27
rect 47 -11 51 -7
rect 118 -11 122 -7
rect 41 -28 45 -24
rect 50 -28 54 -24
rect 66 -47 70 -43
rect 76 -54 80 -50
rect 115 -28 119 -24
rect 99 -47 103 -43
rect 124 -28 128 -24
rect 89 -54 93 -50
<< metal1 >>
rect 35 101 134 104
rect 35 61 38 101
rect 72 71 76 72
rect 83 71 86 98
rect 71 68 86 71
rect 97 68 98 71
rect 35 58 52 61
rect 61 57 65 60
rect 52 52 55 57
rect 71 52 74 68
rect 95 52 98 68
rect 131 61 134 101
rect 104 57 108 60
rect 117 58 134 61
rect 114 52 117 57
rect 52 43 55 48
rect 71 43 74 48
rect 84 42 89 46
rect 95 43 98 48
rect 114 43 117 48
rect 52 34 55 39
rect 35 30 52 33
rect 61 31 65 34
rect 35 -1 38 30
rect 71 23 74 39
rect 95 23 98 39
rect 114 34 117 39
rect 104 31 108 34
rect 117 30 134 33
rect 71 20 86 23
rect 72 19 76 20
rect 83 -1 86 20
rect 97 20 98 23
rect 131 -1 134 30
rect 35 -4 44 -1
rect 41 -14 44 -4
rect 62 -4 86 -1
rect 125 -4 134 -1
rect 55 -11 114 -8
rect 125 -14 128 -4
rect 40 -18 42 -14
rect 54 -18 67 -14
rect 79 -17 90 -14
rect 41 -24 44 -18
rect 51 -24 54 -18
rect 54 -28 56 -24
rect 53 -38 56 -28
rect 64 -27 79 -24
rect 60 -30 63 -27
rect 76 -30 79 -27
rect 39 -45 42 -42
rect 59 -45 62 -34
rect 39 -48 62 -45
rect 59 -54 76 -51
rect 59 -57 62 -54
rect 83 -57 86 -17
rect 102 -18 115 -14
rect 127 -18 129 -14
rect 90 -27 105 -24
rect 115 -24 118 -18
rect 125 -24 128 -18
rect 90 -30 93 -27
rect 106 -30 109 -27
rect 113 -28 115 -24
rect 107 -45 110 -34
rect 113 -38 116 -28
rect 127 -45 130 -42
rect 107 -48 130 -45
rect 93 -54 110 -51
rect 107 -57 110 -54
<< m2contact >>
rect 93 68 97 72
rect 51 64 55 68
rect 45 47 49 51
rect 87 55 91 59
rect 114 64 118 68
rect 45 40 49 44
rect 80 39 84 46
rect 120 47 124 51
rect 51 23 55 27
rect 87 32 91 36
rect 120 40 124 44
rect 114 23 118 27
rect 93 19 97 23
rect 58 -5 62 -1
rect 51 -11 55 -7
rect 114 -11 118 -7
rect 60 -27 64 -23
rect 67 -38 71 -34
rect 70 -47 74 -43
rect 105 -27 109 -23
rect 98 -38 102 -34
rect 95 -47 99 -43
rect 82 -61 86 -57
<< metal2 >>
rect 83 71 86 98
rect 83 68 93 71
rect 19 65 51 68
rect 19 26 22 65
rect 55 65 69 68
rect 100 65 114 68
rect 66 62 103 65
rect 118 65 131 68
rect 29 58 52 61
rect 82 58 87 59
rect 49 55 87 58
rect 117 58 131 61
rect 91 55 120 58
rect 73 49 96 52
rect 73 47 76 49
rect 32 44 76 47
rect 93 47 96 49
rect 93 44 131 47
rect 49 33 87 36
rect 29 30 52 33
rect 82 32 87 33
rect 91 33 120 36
rect 117 30 131 33
rect 19 23 51 26
rect 66 26 103 29
rect 55 23 69 26
rect 100 23 114 26
rect 118 23 131 26
rect 83 20 93 23
rect 83 -1 86 20
rect 62 -5 63 -2
rect 83 -4 109 -1
rect 35 -10 51 -7
rect 47 -11 51 -10
rect 60 -23 63 -5
rect 106 -23 109 -4
rect 118 -10 133 -7
rect 118 -11 122 -10
rect 35 -47 70 -44
rect 74 -47 95 -44
rect 99 -47 133 -44
rect 35 -61 82 -58
rect 86 -61 133 -58
<< m3contact >>
rect 84 39 90 46
rect 71 -39 75 -35
rect 94 -39 98 -35
<< metal3 >>
rect 48 57 70 68
rect 99 57 121 68
rect 48 48 121 57
rect 27 46 142 48
rect 27 43 84 46
rect 27 -34 32 43
rect 48 39 84 43
rect 90 43 142 46
rect 90 39 121 43
rect 48 34 121 39
rect 48 23 70 34
rect 99 23 121 34
rect 137 -34 142 43
rect 27 -35 142 -34
rect 27 -39 71 -35
rect 75 -39 94 -35
rect 98 -39 142 -35
rect 27 -40 142 -39
<< end >>
