magic
tech scmos
timestamp 1354245433
<< ntransistor >>
rect 24 71 27 73
rect 11 64 13 67
rect 66 71 69 73
rect 80 64 82 67
rect 20 54 22 57
rect 30 54 32 57
rect 61 54 63 57
rect 71 54 73 57
rect 20 34 22 37
rect 30 34 32 37
rect 61 34 63 37
rect 71 34 73 37
rect 11 24 13 27
rect 24 18 27 20
rect -103 -26 -100 -24
rect -116 -33 -114 -30
rect 80 24 82 27
rect 66 18 69 20
rect -61 -26 -58 -24
rect -77 -33 -74 -32
rect -47 -33 -45 -30
rect -107 -42 -105 -39
rect -97 -42 -95 -39
rect -66 -42 -64 -39
rect -56 -42 -54 -39
rect -107 -52 -105 -49
rect -97 -52 -95 -49
rect -66 -52 -64 -49
rect -56 -52 -54 -49
rect -116 -61 -114 -58
rect -77 -59 -74 -58
rect -103 -67 -100 -65
rect -47 -61 -45 -58
rect -61 -67 -58 -65
<< ndiffusion >>
rect 0 75 42 92
rect 0 71 16 75
rect 22 74 42 75
rect 0 67 10 71
rect 24 73 27 74
rect 24 70 27 71
rect 0 64 11 67
rect 13 64 14 67
rect 0 62 10 64
rect 0 56 6 62
rect 0 50 10 56
rect 32 62 42 74
rect 51 75 93 92
rect 51 74 71 75
rect 51 62 61 74
rect 66 73 69 74
rect 66 70 69 71
rect 77 71 93 75
rect 83 67 93 71
rect 79 64 80 67
rect 82 64 93 67
rect 18 54 20 57
rect 22 54 30 57
rect 32 54 33 57
rect 83 62 93 64
rect 60 54 61 57
rect 63 54 71 57
rect 73 54 75 57
rect 87 56 93 62
rect 0 35 10 41
rect 83 50 93 56
rect 0 29 6 35
rect 18 34 20 37
rect 22 34 30 37
rect 32 34 33 37
rect 0 27 10 29
rect 60 34 61 37
rect 63 34 71 37
rect 73 34 75 37
rect 0 24 11 27
rect 13 24 14 27
rect 0 20 10 24
rect 0 16 16 20
rect 24 20 27 21
rect 24 17 27 18
rect 32 17 42 29
rect 22 16 42 17
rect -127 -22 -82 1
rect -127 -23 -111 -22
rect -105 -23 -82 -22
rect -127 -30 -117 -23
rect -103 -24 -100 -23
rect -103 -27 -100 -26
rect -127 -33 -116 -30
rect -114 -33 -113 -30
rect -127 -35 -118 -33
rect -127 -41 -121 -35
rect -95 -31 -82 -23
rect -79 -22 -34 1
rect 0 -1 42 16
rect 51 17 61 29
rect 83 35 93 41
rect 87 29 93 35
rect 83 27 93 29
rect 79 24 80 27
rect 82 24 93 27
rect 66 20 69 21
rect 66 17 69 18
rect 83 20 93 24
rect 51 16 71 17
rect 77 16 93 20
rect 51 -1 93 16
rect -79 -23 -56 -22
rect -50 -23 -34 -22
rect -79 -31 -66 -23
rect -61 -24 -58 -23
rect -61 -27 -58 -26
rect -44 -30 -34 -23
rect -95 -33 -84 -31
rect -77 -32 -66 -31
rect -74 -33 -66 -32
rect -48 -33 -47 -30
rect -45 -33 -34 -30
rect -43 -35 -34 -33
rect -127 -44 -117 -41
rect -109 -42 -107 -39
rect -105 -42 -97 -39
rect -95 -42 -94 -39
rect -67 -42 -66 -39
rect -64 -42 -56 -39
rect -54 -42 -52 -39
rect -40 -41 -34 -35
rect -44 -44 -34 -41
rect -127 -50 -117 -47
rect -127 -56 -121 -50
rect -109 -52 -107 -49
rect -105 -52 -97 -49
rect -95 -52 -94 -49
rect -127 -58 -118 -56
rect -67 -52 -66 -49
rect -64 -52 -56 -49
rect -54 -52 -52 -49
rect -44 -50 -34 -47
rect -127 -61 -116 -58
rect -114 -61 -113 -58
rect -95 -60 -84 -58
rect -74 -59 -66 -58
rect -77 -60 -66 -59
rect -127 -68 -117 -61
rect -103 -65 -100 -64
rect -103 -68 -100 -67
rect -95 -68 -82 -60
rect -127 -69 -111 -68
rect -105 -69 -82 -68
rect -127 -92 -82 -69
rect -79 -68 -66 -60
rect -40 -56 -34 -50
rect -43 -58 -34 -56
rect -48 -61 -47 -58
rect -45 -61 -34 -58
rect -61 -65 -58 -64
rect -61 -68 -58 -67
rect -44 -68 -34 -61
rect -79 -69 -56 -68
rect -50 -69 -34 -68
rect -79 -92 -34 -69
<< ndcontact >>
rect 14 63 18 67
rect 24 66 28 70
rect 14 54 18 58
rect 65 66 69 70
rect 75 63 79 67
rect 33 54 37 58
rect 56 54 60 58
rect 75 54 79 58
rect 14 33 18 37
rect 33 33 37 37
rect 56 33 60 37
rect 14 24 18 28
rect 24 21 28 25
rect -113 -34 -109 -30
rect -103 -31 -99 -27
rect 75 33 79 37
rect 65 21 69 25
rect 75 24 79 28
rect -62 -31 -58 -27
rect -52 -34 -48 -30
rect -113 -43 -109 -39
rect -94 -43 -90 -39
rect -71 -43 -67 -39
rect -52 -43 -48 -39
rect -113 -52 -109 -48
rect -94 -52 -90 -48
rect -71 -52 -67 -48
rect -52 -52 -48 -48
rect -113 -61 -109 -57
rect -103 -64 -99 -60
rect -62 -64 -58 -60
rect -52 -61 -48 -57
<< psubstratepdiff >>
rect 38 49 55 50
rect 38 42 39 49
rect 43 42 55 49
rect 38 41 55 42
rect -86 -39 -75 -37
rect -86 -45 -85 -39
rect -76 -45 -75 -39
rect -86 -54 -75 -45
<< psubstratepcontact >>
rect 39 42 43 49
rect -85 -45 -76 -39
<< polysilicon >>
rect 21 71 24 73
rect 27 71 29 73
rect 11 67 13 69
rect 11 58 13 64
rect 20 57 22 61
rect 64 71 66 73
rect 69 71 72 73
rect 80 67 82 69
rect 30 57 32 59
rect 61 57 63 59
rect 71 57 73 61
rect 80 58 82 64
rect 20 52 22 54
rect 30 49 32 54
rect 61 49 63 54
rect 71 52 73 54
rect 20 37 22 39
rect 30 37 32 42
rect 61 37 63 42
rect 71 37 73 39
rect 11 27 13 33
rect 20 30 22 34
rect 30 32 32 34
rect 61 32 63 34
rect 11 22 13 24
rect 21 18 24 20
rect 27 18 29 20
rect -106 -26 -103 -24
rect -100 -26 -98 -24
rect -116 -30 -114 -28
rect -116 -39 -114 -33
rect 71 30 73 34
rect 80 27 82 33
rect 80 22 82 24
rect 64 18 66 20
rect 69 18 72 20
rect -63 -26 -61 -24
rect -58 -26 -55 -24
rect -47 -30 -45 -28
rect -107 -39 -105 -36
rect -97 -36 -83 -34
rect -78 -33 -77 -32
rect -78 -34 -74 -33
rect -78 -36 -64 -34
rect -97 -39 -95 -36
rect -66 -39 -64 -36
rect -56 -39 -54 -36
rect -47 -39 -45 -33
rect -107 -44 -105 -42
rect -97 -44 -95 -42
rect -66 -44 -64 -42
rect -56 -44 -54 -42
rect -107 -49 -105 -47
rect -97 -49 -95 -47
rect -116 -58 -114 -52
rect -107 -55 -105 -52
rect -97 -55 -95 -52
rect -66 -49 -64 -47
rect -56 -49 -54 -47
rect -66 -55 -64 -52
rect -97 -57 -83 -55
rect -78 -57 -64 -55
rect -56 -55 -54 -52
rect -78 -58 -74 -57
rect -78 -59 -77 -58
rect -116 -63 -114 -61
rect -106 -67 -103 -65
rect -100 -67 -98 -65
rect -47 -58 -45 -52
rect -47 -63 -45 -61
rect -63 -67 -61 -65
rect -58 -67 -55 -65
<< polycontact >>
rect 17 70 21 74
rect 7 57 11 61
rect 22 59 26 63
rect 72 70 76 74
rect 67 59 71 63
rect 82 57 86 61
rect 26 48 30 52
rect 26 39 30 43
rect 63 48 67 52
rect 63 39 67 43
rect 7 30 11 34
rect 22 28 26 32
rect 17 17 21 21
rect -110 -27 -106 -23
rect -120 -40 -116 -36
rect 67 28 71 32
rect 82 30 86 34
rect 72 17 76 21
rect -55 -27 -51 -23
rect -105 -38 -101 -34
rect -83 -36 -78 -32
rect -60 -38 -56 -34
rect -45 -40 -41 -36
rect -120 -55 -116 -51
rect -105 -57 -101 -53
rect -83 -59 -78 -55
rect -60 -57 -56 -53
rect -110 -68 -106 -64
rect -45 -55 -41 -51
rect -55 -68 -51 -64
<< metal1 >>
rect 7 67 10 92
rect 7 64 14 67
rect 23 63 27 66
rect 14 58 17 63
rect 42 58 45 92
rect 37 55 45 58
rect 48 58 51 92
rect 83 67 86 92
rect 66 63 70 66
rect 79 64 86 67
rect 76 58 79 63
rect 48 55 56 58
rect 14 50 17 54
rect 7 47 17 50
rect 33 47 36 54
rect 7 41 17 44
rect 14 37 17 41
rect 33 37 36 44
rect 57 47 60 54
rect 76 50 79 54
rect 76 47 86 50
rect 57 37 60 44
rect 76 41 86 44
rect 76 37 79 41
rect 37 33 45 36
rect 14 28 17 33
rect 7 24 14 27
rect 23 25 27 28
rect -130 -30 -127 4
rect -130 -33 -113 -30
rect -104 -34 -100 -31
rect -113 -39 -110 -34
rect -94 -39 -91 4
rect -70 -39 -67 4
rect 7 -1 10 24
rect 42 -1 45 33
rect 48 33 56 36
rect 48 -1 51 33
rect 76 28 79 33
rect 66 25 70 28
rect 79 24 86 27
rect 83 -1 86 24
rect -61 -34 -57 -31
rect -48 -33 -34 -30
rect -51 -39 -48 -34
rect -113 -48 -110 -43
rect -94 -48 -91 -43
rect -81 -49 -76 -45
rect -70 -48 -67 -43
rect -51 -48 -48 -43
rect -113 -57 -110 -52
rect -130 -61 -113 -58
rect -104 -60 -100 -57
rect -130 -92 -127 -61
rect -94 -92 -91 -52
rect -70 -92 -67 -52
rect -51 -57 -48 -52
rect -61 -60 -57 -57
rect -48 -61 -34 -58
<< m2contact >>
rect 13 70 17 74
rect 7 53 11 57
rect 76 70 80 74
rect 22 47 26 51
rect 7 34 11 38
rect 22 40 26 44
rect 43 43 47 48
rect 67 47 71 51
rect 82 53 86 57
rect 67 40 71 44
rect -114 -27 -110 -23
rect -120 -44 -116 -40
rect -78 -36 -74 -32
rect 13 17 17 21
rect 82 34 86 38
rect 76 17 80 21
rect -51 -27 -47 -23
rect -120 -51 -116 -47
rect -85 -52 -81 -45
rect -45 -44 -41 -40
rect -114 -68 -110 -64
rect -78 -59 -74 -55
rect -45 -51 -41 -47
rect -51 -68 -47 -64
<< metal2 >>
rect 0 71 13 74
rect 17 71 45 74
rect 48 71 76 74
rect 80 71 93 74
rect 0 57 45 60
rect 48 57 93 60
rect 22 51 45 54
rect 48 51 71 54
rect 0 47 22 50
rect 0 41 22 44
rect 71 47 93 50
rect 71 41 93 44
rect 22 37 45 40
rect 48 37 71 40
rect 0 31 45 34
rect 48 31 93 34
rect 0 17 13 20
rect 17 17 45 20
rect 48 17 76 20
rect 80 17 93 20
rect -130 -26 -114 -23
rect -110 -26 -51 -23
rect -47 -26 -34 -23
rect -83 -33 -78 -32
rect -130 -36 -78 -33
rect -74 -36 -34 -33
rect -92 -42 -69 -39
rect -92 -44 -89 -42
rect -130 -47 -89 -44
rect -72 -44 -69 -42
rect -72 -47 -34 -44
rect -130 -58 -78 -55
rect -83 -59 -78 -58
rect -74 -58 -34 -55
rect -130 -68 -114 -65
rect -110 -68 -51 -65
rect -47 -68 -34 -65
<< m3contact >>
rect 47 43 51 48
rect -81 -52 -75 -45
<< metal3 >>
rect 46 48 52 49
rect 46 43 47 48
rect 51 43 52 48
rect 46 42 52 43
rect -117 -34 -95 -23
rect -66 -34 -44 -23
rect -117 -43 -44 -34
rect -130 -45 -34 -43
rect -130 -48 -81 -45
rect -117 -52 -81 -48
rect -75 -48 -34 -45
rect -75 -52 -44 -48
rect -117 -57 -44 -52
rect -117 -68 -95 -57
rect -66 -68 -44 -57
<< labels >>
rlabel metal1 50 91 50 91 5 Column
rlabel metal1 85 91 85 91 5 Vdd
rlabel metal2 49 52 49 52 1 Row
rlabel metal2 92 58 92 58 7 Reset
rlabel metal2 92 72 92 72 7 Shutter
rlabel metal2 -35 -25 -35 -25 7 Shutter
rlabel metal2 -36 -35 -36 -35 1 Row
rlabel metal2 -37 -45 -37 -45 1 Reset
rlabel metal1 -69 -3 -69 -3 1 Column
rlabel metal2 -126 -25 -126 -25 3 Shutter
rlabel metal2 -125 -35 -125 -35 1 Row
rlabel metal2 -124 -45 -124 -45 1 Reset
rlabel metal1 -92 -3 -92 -3 1 Column
rlabel metal1 -128 -3 -128 -3 1 Vdd
rlabel metal2 -35 -66 -35 -66 7 Shutter
rlabel metal2 -36 -56 -36 -56 5 Row
rlabel metal2 -37 -46 -37 -46 5 Reset
rlabel metal1 -69 -88 -69 -88 5 Column
rlabel metal2 -126 -66 -126 -66 3 Shutter
rlabel metal2 -125 -56 -125 -56 5 Row
rlabel metal2 -124 -46 -124 -46 5 Reset
rlabel metal1 -92 -88 -92 -88 5 Column
rlabel metal1 -128 -88 -128 -88 5 Vdd
<< end >>
