magic
tech scmos
timestamp 1355369891
<< nwell >>
rect -69 2979 -20 3101
<< pwell >>
rect -116 2979 -69 3101
<< ntransistor >>
rect -103 3050 -97 3058
rect -81 3050 -75 3058
rect -103 3042 -97 3044
rect -81 3042 -75 3044
rect -103 3034 -97 3036
rect -81 3034 -75 3036
rect -103 3029 -97 3031
rect -81 3029 -75 3031
rect -103 3013 -97 3021
rect -81 3013 -75 3021
rect -103 3005 -97 3007
rect -81 3005 -75 3007
rect -103 2997 -97 2999
rect -81 2997 -75 2999
rect -103 2992 -97 2994
rect -81 2992 -75 2994
<< ptransistor >>
rect -63 3056 -57 3058
rect -41 3056 -35 3058
rect -63 3051 -57 3053
rect -41 3051 -35 3053
rect -63 3037 -57 3045
rect -41 3037 -35 3045
rect -63 3029 -57 3031
rect -41 3029 -35 3031
rect -63 3019 -57 3021
rect -41 3019 -35 3021
rect -63 3014 -57 3016
rect -41 3014 -35 3016
rect -63 3000 -57 3008
rect -41 3000 -35 3008
rect -63 2992 -57 2994
rect -41 2992 -35 2994
<< ndiffusion >>
rect -103 3058 -97 3095
rect -81 3058 -75 3095
rect -103 3049 -97 3050
rect -103 3045 -102 3049
rect -98 3045 -97 3049
rect -103 3044 -97 3045
rect -81 3049 -75 3050
rect -81 3045 -80 3049
rect -76 3045 -75 3049
rect -81 3044 -75 3045
rect -103 3041 -97 3042
rect -103 3037 -102 3041
rect -98 3037 -97 3041
rect -81 3041 -75 3042
rect -81 3037 -80 3041
rect -76 3037 -75 3041
rect -103 3036 -97 3037
rect -81 3036 -75 3037
rect -103 3031 -97 3034
rect -81 3031 -75 3034
rect -103 3028 -97 3029
rect -103 3024 -102 3028
rect -98 3024 -97 3028
rect -103 3021 -97 3024
rect -81 3028 -75 3029
rect -81 3024 -80 3028
rect -76 3024 -75 3028
rect -81 3021 -75 3024
rect -103 3012 -97 3013
rect -103 3008 -102 3012
rect -98 3008 -97 3012
rect -103 3007 -97 3008
rect -81 3012 -75 3013
rect -81 3008 -80 3012
rect -76 3008 -75 3012
rect -81 3007 -75 3008
rect -103 3004 -97 3005
rect -103 3000 -102 3004
rect -98 3000 -97 3004
rect -81 3004 -75 3005
rect -81 3000 -80 3004
rect -76 3000 -75 3004
rect -103 2999 -97 3000
rect -81 2999 -75 3000
rect -103 2994 -97 2997
rect -81 2994 -75 2997
rect -103 2991 -97 2992
rect -103 2987 -102 2991
rect -98 2987 -97 2991
rect -103 2985 -97 2987
rect -81 2991 -75 2992
rect -81 2987 -80 2991
rect -76 2987 -75 2991
rect -81 2985 -75 2987
<< pdiffusion >>
rect -63 3058 -57 3095
rect -41 3058 -35 3095
rect -63 3053 -57 3056
rect -41 3053 -35 3056
rect -63 3050 -57 3051
rect -63 3046 -62 3050
rect -58 3046 -57 3050
rect -63 3045 -57 3046
rect -41 3050 -35 3051
rect -41 3046 -40 3050
rect -36 3046 -35 3050
rect -41 3045 -35 3046
rect -63 3036 -57 3037
rect -63 3032 -62 3036
rect -58 3032 -57 3036
rect -63 3031 -57 3032
rect -41 3036 -35 3037
rect -41 3032 -40 3036
rect -36 3032 -35 3036
rect -41 3031 -35 3032
rect -63 3028 -57 3029
rect -63 3024 -62 3028
rect -58 3024 -57 3028
rect -41 3028 -35 3029
rect -41 3024 -40 3028
rect -36 3024 -35 3028
rect -63 3021 -57 3024
rect -41 3021 -35 3024
rect -63 3016 -57 3019
rect -41 3016 -35 3019
rect -63 3013 -57 3014
rect -63 3009 -62 3013
rect -58 3009 -57 3013
rect -63 3008 -57 3009
rect -41 3013 -35 3014
rect -41 3009 -40 3013
rect -36 3009 -35 3013
rect -41 3008 -35 3009
rect -63 2999 -57 3000
rect -63 2995 -62 2999
rect -58 2995 -57 2999
rect -63 2994 -57 2995
rect -41 2999 -35 3000
rect -41 2995 -40 2999
rect -36 2995 -35 2999
rect -41 2994 -35 2995
rect -63 2991 -57 2992
rect -63 2987 -62 2991
rect -58 2987 -57 2991
rect -41 2991 -35 2992
rect -41 2987 -40 2991
rect -36 2987 -35 2991
rect -63 2985 -57 2987
rect -41 2985 -35 2987
<< ndcontact >>
rect -102 3045 -98 3049
rect -80 3045 -76 3049
rect -102 3037 -98 3041
rect -80 3037 -76 3041
rect -102 3024 -98 3028
rect -80 3024 -76 3028
rect -102 3008 -98 3012
rect -80 3008 -76 3012
rect -102 3000 -98 3004
rect -80 3000 -76 3004
rect -102 2987 -98 2991
rect -80 2987 -76 2991
<< pdcontact >>
rect -62 3046 -58 3050
rect -40 3046 -36 3050
rect -62 3032 -58 3036
rect -40 3032 -36 3036
rect -62 3024 -58 3028
rect -40 3024 -36 3028
rect -62 3009 -58 3013
rect -40 3009 -36 3013
rect -62 2995 -58 2999
rect -40 2995 -36 2999
rect -62 2987 -58 2991
rect -40 2987 -36 2991
<< psubstratepdiff >>
rect -92 3042 -86 3043
rect -92 3038 -91 3042
rect -87 3038 -86 3042
rect -92 3037 -86 3038
rect -92 3005 -86 3006
rect -92 3001 -91 3005
rect -87 3001 -86 3005
rect -92 3000 -86 3001
<< nsubstratendiff >>
rect -52 3029 -46 3030
rect -52 3025 -51 3029
rect -47 3025 -46 3029
rect -52 3024 -46 3025
rect -52 2992 -46 2993
rect -52 2988 -51 2992
rect -47 2988 -46 2992
rect -52 2987 -46 2988
<< psubstratepcontact >>
rect -91 3038 -87 3042
rect -91 3001 -87 3005
<< nsubstratencontact >>
rect -51 3025 -47 3029
rect -51 2988 -47 2992
<< polysilicon >>
rect -116 3055 -110 3056
rect -105 3055 -103 3058
rect -116 3051 -115 3055
rect -111 3053 -103 3055
rect -111 3051 -110 3053
rect -116 3050 -110 3051
rect -105 3050 -103 3053
rect -97 3055 -95 3058
rect -83 3055 -81 3058
rect -97 3053 -81 3055
rect -97 3050 -95 3053
rect -83 3050 -81 3053
rect -75 3056 -63 3058
rect -57 3056 -41 3058
rect -35 3056 -33 3058
rect -30 3056 -24 3057
rect -75 3050 -73 3056
rect -30 3053 -29 3056
rect -70 3051 -63 3053
rect -57 3051 -50 3053
rect -43 3051 -41 3053
rect -35 3052 -29 3053
rect -25 3052 -24 3056
rect -35 3051 -24 3052
rect -115 3036 -113 3050
rect -110 3044 -104 3045
rect -92 3049 -86 3050
rect -92 3045 -91 3049
rect -87 3046 -86 3049
rect -87 3045 -82 3046
rect -92 3044 -82 3045
rect -70 3044 -68 3051
rect -52 3050 -46 3051
rect -52 3046 -51 3050
rect -47 3046 -46 3050
rect -52 3045 -46 3046
rect -110 3040 -109 3044
rect -105 3042 -103 3044
rect -97 3042 -95 3044
rect -84 3042 -81 3044
rect -75 3042 -68 3044
rect -105 3040 -104 3042
rect -110 3039 -104 3040
rect -65 3039 -63 3045
rect -70 3037 -63 3039
rect -57 3042 -55 3045
rect -43 3042 -41 3045
rect -57 3040 -41 3042
rect -57 3037 -55 3040
rect -43 3037 -41 3040
rect -35 3037 -33 3045
rect -70 3036 -68 3037
rect -115 3034 -103 3036
rect -97 3034 -81 3036
rect -75 3034 -68 3036
rect -52 3036 -46 3037
rect -52 3033 -51 3036
rect -56 3032 -51 3033
rect -47 3032 -46 3036
rect -56 3031 -46 3032
rect -30 3034 -24 3035
rect -30 3031 -29 3034
rect -114 3030 -103 3031
rect -114 3026 -113 3030
rect -109 3029 -103 3030
rect -97 3029 -95 3031
rect -88 3029 -81 3031
rect -75 3029 -63 3031
rect -57 3029 -54 3031
rect -43 3029 -41 3031
rect -35 3030 -29 3031
rect -25 3030 -24 3034
rect -35 3029 -24 3030
rect -109 3026 -108 3029
rect -114 3025 -108 3026
rect -92 3028 -86 3029
rect -92 3024 -91 3028
rect -87 3024 -86 3028
rect -92 3023 -86 3024
rect -116 3018 -110 3019
rect -105 3018 -103 3021
rect -116 3014 -115 3018
rect -111 3016 -103 3018
rect -111 3014 -110 3016
rect -116 3013 -110 3014
rect -105 3013 -103 3016
rect -97 3018 -95 3021
rect -83 3018 -81 3021
rect -97 3016 -81 3018
rect -97 3013 -95 3016
rect -83 3013 -81 3016
rect -75 3019 -63 3021
rect -57 3019 -41 3021
rect -35 3019 -33 3021
rect -30 3019 -24 3020
rect -75 3013 -73 3019
rect -30 3016 -29 3019
rect -70 3014 -63 3016
rect -57 3014 -50 3016
rect -43 3014 -41 3016
rect -35 3015 -29 3016
rect -25 3015 -24 3019
rect -35 3014 -24 3015
rect -115 2999 -113 3013
rect -110 3007 -104 3008
rect -92 3012 -86 3013
rect -92 3008 -91 3012
rect -87 3009 -86 3012
rect -87 3008 -82 3009
rect -92 3007 -82 3008
rect -70 3007 -68 3014
rect -52 3013 -46 3014
rect -52 3009 -51 3013
rect -47 3009 -46 3013
rect -52 3008 -46 3009
rect -110 3003 -109 3007
rect -105 3005 -103 3007
rect -97 3005 -95 3007
rect -84 3005 -81 3007
rect -75 3005 -68 3007
rect -105 3003 -104 3005
rect -110 3002 -104 3003
rect -65 3002 -63 3008
rect -70 3000 -63 3002
rect -57 3005 -55 3008
rect -43 3005 -41 3008
rect -57 3003 -41 3005
rect -57 3000 -55 3003
rect -43 3000 -41 3003
rect -35 3000 -33 3008
rect -70 2999 -68 3000
rect -115 2997 -103 2999
rect -97 2997 -81 2999
rect -75 2997 -68 2999
rect -52 2999 -46 3000
rect -52 2996 -51 2999
rect -56 2995 -51 2996
rect -47 2995 -46 2999
rect -56 2994 -46 2995
rect -30 2997 -24 2998
rect -30 2994 -29 2997
rect -114 2993 -103 2994
rect -114 2989 -113 2993
rect -109 2992 -103 2993
rect -97 2992 -95 2994
rect -88 2992 -81 2994
rect -75 2992 -63 2994
rect -57 2992 -54 2994
rect -43 2992 -41 2994
rect -35 2993 -29 2994
rect -25 2993 -24 2997
rect -35 2992 -24 2993
rect -109 2989 -108 2992
rect -114 2988 -108 2989
rect -92 2991 -86 2992
rect -92 2987 -91 2991
rect -87 2987 -86 2991
rect -92 2986 -86 2987
<< polycontact >>
rect -115 3051 -111 3055
rect -29 3052 -25 3056
rect -91 3045 -87 3049
rect -51 3046 -47 3050
rect -109 3040 -105 3044
rect -51 3032 -47 3036
rect -113 3026 -109 3030
rect -29 3030 -25 3034
rect -91 3024 -87 3028
rect -115 3014 -111 3018
rect -29 3015 -25 3019
rect -91 3008 -87 3012
rect -51 3009 -47 3013
rect -109 3003 -105 3007
rect -51 2995 -47 2999
rect -113 2989 -109 2993
rect -29 2993 -25 2997
rect -91 2987 -87 2991
<< metal1 >>
rect -108 3053 -29 3056
rect -108 3044 -105 3053
rect -80 3049 -76 3053
rect -98 3045 -91 3049
rect -62 3050 -58 3053
rect -47 3046 -40 3050
rect -98 3037 -97 3041
rect -93 3038 -91 3041
rect -87 3038 -85 3041
rect -93 3037 -85 3038
rect -81 3037 -80 3041
rect -62 3039 -20 3043
rect -62 3036 -58 3039
rect -112 3032 -62 3034
rect -47 3032 -40 3036
rect -29 3034 -26 3039
rect -112 3031 -58 3032
rect -112 3030 -109 3031
rect -80 3028 -76 3031
rect -98 3024 -91 3028
rect -58 3024 -57 3028
rect -53 3025 -51 3028
rect -47 3025 -45 3028
rect -53 3024 -45 3025
rect -41 3024 -40 3028
rect -13 3025 -10 3095
rect -108 3016 -29 3019
rect -108 3007 -105 3016
rect -80 3012 -76 3016
rect -98 3008 -91 3012
rect -62 3013 -58 3016
rect -47 3009 -40 3013
rect -98 3000 -97 3004
rect -93 3001 -91 3004
rect -87 3001 -85 3004
rect -93 3000 -85 3001
rect -81 3000 -80 3004
rect -62 3002 -20 3006
rect -62 2999 -58 3002
rect -112 2995 -62 2997
rect -47 2995 -40 2999
rect -29 2997 -26 3002
rect -112 2994 -58 2995
rect -112 2993 -109 2994
rect -80 2991 -76 2994
rect -98 2987 -91 2991
rect -58 2987 -57 2991
rect -53 2988 -51 2991
rect -47 2988 -45 2991
rect -53 2987 -45 2988
rect -41 2987 -40 2991
rect -13 2987 -10 3021
rect -7 3045 -4 3095
rect -7 3004 -4 3041
rect -7 2987 -4 3000
<< m2contact >>
rect -115 3047 -111 3051
rect -97 3037 -93 3041
rect -85 3037 -81 3041
rect -20 3038 -16 3042
rect -57 3024 -53 3028
rect -45 3024 -41 3028
rect -14 3021 -10 3025
rect -115 3010 -111 3014
rect -97 3000 -93 3004
rect -85 3000 -81 3004
rect -20 3003 -16 3007
rect -57 2987 -53 2991
rect -45 2987 -41 2991
rect -7 3041 -3 3045
rect -7 3000 -3 3004
<< metal2 >>
rect -115 3051 -111 3101
rect -115 3014 -111 3047
rect -115 2985 -111 3010
rect -98 3041 -80 3101
rect -98 3037 -97 3041
rect -93 3037 -85 3041
rect -81 3037 -80 3041
rect -98 3004 -80 3037
rect -98 3000 -97 3004
rect -93 3000 -85 3004
rect -81 3000 -80 3004
rect -98 2985 -80 3000
rect -58 3028 -40 3101
rect -20 3034 -3 3038
rect -58 3024 -57 3028
rect -53 3024 -45 3028
rect -41 3024 -40 3028
rect -58 2991 -40 3024
rect -10 3021 -3 3024
rect -20 3007 -3 3011
rect -58 2987 -57 2991
rect -53 2987 -45 2991
rect -41 2987 -40 2991
rect -58 2985 -40 2987
<< metal3 >>
rect -20 3025 -4 3101
rect -20 3020 -3 3025
rect -20 2987 -4 3020
<< labels >>
rlabel pdiffusion -38 3060 -38 3060 5 pos1
rlabel pdiffusion -60 3060 -60 3060 5 pos2
rlabel metal2 -45 3030 -45 3030 3 pos
rlabel metal2 -89 3057 -89 3057 5 neg
rlabel ndiffusion -78 3060 -78 3060 5 d
rlabel ndiffusion -100 3060 -100 3060 5 db
rlabel ndcontact -78 3025 -78 3025 1 q
rlabel ndcontact -100 3025 -100 3025 1 qb
rlabel ndiffusion -100 3024 -100 3024 5 db
rlabel ndiffusion -78 3024 -78 3024 5 d
rlabel pdiffusion -60 3024 -60 3024 5 pos2
rlabel pdiffusion -38 3024 -38 3024 5 pos1
rlabel metal2 -113 3024 -113 3024 2 clk
rlabel metal2 -113 2987 -113 2987 2 clk
rlabel ndcontact -100 2988 -100 2988 1 qb
rlabel ndcontact -78 2988 -78 2988 1 q
rlabel metal2 -89 3020 -89 3020 5 neg
rlabel metal2 -45 2993 -45 2993 3 pos
rlabel metal3 -18 3093 -18 3093 1 Gnd
rlabel metal1 -6 3094 -6 3094 5 Shutter
rlabel metal1 -11 3094 -11 3094 5 Reset
<< end >>
