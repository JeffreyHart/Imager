magic
tech scmos
timestamp 1355375890
<< polysilicon >>
rect 4295 602 4298 604
rect 4293 573 4298 575
<< polycontact >>
rect 4291 602 4295 606
rect 4289 573 4293 577
<< metal1 >>
rect 1013 4359 1053 4487
rect 671 4346 1053 4359
rect 704 4322 720 4325
rect 1013 4318 1053 4346
rect 1487 4318 1527 4487
rect 1961 4318 2001 4487
rect 2435 4318 2475 4487
rect 2909 4318 2949 4487
rect 3383 4318 3423 4487
rect 3857 4318 3897 4487
rect 711 4308 4266 4318
rect 711 4302 714 4308
rect 759 4302 762 4308
rect 807 4302 810 4308
rect 855 4302 858 4308
rect 903 4302 906 4308
rect 951 4302 954 4308
rect 999 4302 1002 4308
rect 1047 4302 1050 4308
rect 1095 4302 1098 4308
rect 1143 4302 1146 4308
rect 1191 4302 1194 4308
rect 1239 4302 1242 4308
rect 1287 4302 1290 4308
rect 1335 4302 1338 4308
rect 1383 4302 1386 4308
rect 1431 4302 1434 4308
rect 1479 4302 1482 4308
rect 1527 4302 1530 4308
rect 1575 4302 1578 4308
rect 1623 4302 1626 4308
rect 1671 4302 1674 4308
rect 1719 4302 1722 4308
rect 1767 4302 1770 4308
rect 1815 4302 1818 4308
rect 1863 4302 1866 4308
rect 1911 4302 1914 4308
rect 1959 4302 1962 4308
rect 2007 4302 2010 4308
rect 2055 4302 2058 4308
rect 2103 4302 2106 4308
rect 2151 4302 2154 4308
rect 2199 4302 2202 4308
rect 2247 4302 2250 4308
rect 2295 4302 2298 4308
rect 2343 4302 2346 4308
rect 2391 4302 2394 4308
rect 2439 4302 2442 4308
rect 2487 4302 2490 4308
rect 2535 4302 2538 4308
rect 2583 4302 2586 4308
rect 2631 4302 2634 4308
rect 2679 4302 2682 4308
rect 2727 4302 2730 4308
rect 2775 4302 2778 4308
rect 2823 4302 2826 4308
rect 2871 4302 2874 4308
rect 2919 4302 2922 4308
rect 2967 4302 2970 4308
rect 3015 4302 3018 4308
rect 3063 4302 3066 4308
rect 3111 4302 3114 4308
rect 3159 4302 3162 4308
rect 3207 4302 3210 4308
rect 3255 4302 3258 4308
rect 3303 4302 3306 4308
rect 3351 4302 3354 4308
rect 3399 4302 3402 4308
rect 3447 4302 3450 4308
rect 3495 4302 3498 4308
rect 3543 4302 3546 4308
rect 3591 4302 3594 4308
rect 3639 4302 3642 4308
rect 3687 4302 3690 4308
rect 3735 4302 3738 4308
rect 3783 4302 3786 4308
rect 3831 4302 3834 4308
rect 3879 4302 3882 4308
rect 3927 4302 3930 4308
rect 3975 4302 3978 4308
rect 4023 4302 4026 4308
rect 4071 4302 4074 4308
rect 4119 4302 4122 4308
rect 4167 4302 4170 4308
rect 4215 4302 4218 4308
rect 4263 4302 4266 4308
rect 513 1070 565 1086
rect 559 747 565 1070
rect 631 747 635 758
rect 559 741 635 747
rect 676 735 687 741
rect 521 729 682 735
rect 521 669 527 729
rect 513 629 527 669
rect 4251 524 4255 599
rect 4274 577 4278 686
rect 4291 619 4487 625
rect 4291 606 4295 619
rect 4274 573 4289 577
rect 4251 520 4404 524
rect 4388 513 4404 520
<< m2contact >>
rect 653 4346 671 4359
rect 695 4322 701 4328
rect 720 4322 726 4328
rect 4274 686 4278 690
rect 4359 611 4366 615
<< metal2 >>
rect 595 4454 612 4489
rect 595 4445 640 4454
rect 1071 4451 1086 4487
rect 636 4346 640 4445
rect 695 4445 1086 4451
rect 695 4328 701 4445
rect 1544 4422 1560 4487
rect 720 4416 1560 4422
rect 720 4328 726 4416
rect 513 1544 596 1560
rect 536 710 687 719
rect 536 612 545 710
rect 4264 687 4274 690
rect 4264 666 4360 671
rect 4264 653 4487 666
rect 513 596 545 612
rect 647 636 682 640
rect 647 524 653 636
rect 4359 629 4487 653
rect 4359 615 4366 629
rect 4382 614 4481 619
rect 4474 612 4481 614
rect 4474 596 4491 612
rect 596 518 653 524
rect 596 513 612 518
rect 1070 513 1086 596
<< m3contact >>
rect 673 4471 713 4487
rect 613 4346 631 4359
rect 658 613 682 631
<< metal3 >>
rect 593 4487 714 4488
rect 593 4471 673 4487
rect 713 4471 714 4487
rect 593 4359 714 4471
rect 593 4346 613 4359
rect 631 4346 714 4359
rect 593 740 714 4346
rect 593 631 4313 740
rect 593 613 658 631
rect 682 613 4313 631
rect 593 608 4313 613
rect 593 584 4471 608
rect 4290 537 4471 584
use inpad  inpad_3
timestamp 1259953556
transform -1 0 841 0 -1 5000
box -2 0 476 513
use inpad  inpad_4
timestamp 1259953556
transform -1 0 1315 0 -1 5000
box -2 0 476 513
use inpad  inpad_5
timestamp 1259953556
transform -1 0 1789 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_14
timestamp 1259953556
transform -1 0 2263 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_15
timestamp 1259953556
transform -1 0 2737 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_16
timestamp 1259953556
transform -1 0 3211 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_17
timestamp 1259953556
transform -1 0 3685 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_10
timestamp 1259953556
transform -1 0 4159 0 -1 5000
box -2 0 476 513
use blankpad  blankpad_9
timestamp 1259953556
transform -1 0 4633 0 -1 5000
box -2 0 476 513
use padframe_top  padframe_top_0
timestamp 1259953556
transform 1 0 0 0 1 4487
box 0 0 5000 513
use blankpad  blankpad_27
timestamp 1259953556
transform 0 1 0 -1 0 4633
box -2 0 476 513
use blankpad  blankpad_28
timestamp 1259953556
transform 0 1 0 -1 0 4159
box -2 0 476 513
use blankpad  blankpad_35
timestamp 1259953556
transform 0 1 0 -1 0 3685
box -2 0 476 513
use blankpad  blankpad_34
timestamp 1259953556
transform 0 1 0 -1 0 3211
box -2 0 476 513
use blankpad  blankpad_33
timestamp 1259953556
transform 0 1 0 -1 0 2737
box -2 0 476 513
use blankpad  blankpad_32
timestamp 1259953556
transform 0 1 0 -1 0 2263
box -2 0 476 513
use inorpad  inorpad_3
timestamp 1259953556
transform 0 1 0 -1 0 1789
box -2 0 476 513
use inorpad  inorpad_2
timestamp 1259953556
transform 0 1 0 -1 0 1315
box -2 0 476 513
use imager_nopads  imager_nopads_0
timestamp 1355375323
transform 1 0 711 0 1 747
box -116 -152 3558 3599
use blankpad  blankpad_2
timestamp 1259953556
transform 0 -1 5000 1 0 4159
box -2 0 476 513
use blankpad  blankpad_3
timestamp 1259953556
transform 0 -1 5000 1 0 3685
box -2 0 476 513
use blankpad  blankpad_4
timestamp 1259953556
transform 0 -1 5000 1 0 3211
box -2 0 476 513
use blankpad  blankpad_5
timestamp 1259953556
transform 0 -1 5000 1 0 2737
box -2 0 476 513
use blankpad  blankpad_6
timestamp 1259953556
transform 0 -1 5000 1 0 2263
box -2 0 476 513
use blankpad  blankpad_7
timestamp 1259953556
transform 0 -1 5000 1 0 1789
box -2 0 476 513
use blankpad  blankpad_8
timestamp 1259953556
transform 0 -1 5000 1 0 1315
box -2 0 476 513
use blankpad  blankpad_1
timestamp 1259953556
transform 0 -1 5000 1 0 841
box -2 0 476 513
use diffamp  diffamp_0
timestamp 1355272872
transform 1 0 4318 0 1 486
box -20 51 152 128
use padframe_left  padframe_left_0
timestamp 1259953556
transform 1 0 0 0 1 367
box 2 2 513 4264
use inpad  inpad_2
timestamp 1259953556
transform 0 1 0 -1 0 841
box -2 0 476 513
use inpad  inpad_1
timestamp 1259953556
transform 1 0 367 0 1 0
box -2 0 476 513
use inpad  inpad_0
timestamp 1259953556
transform 1 0 841 0 1 0
box -2 0 476 513
use blankpad  blankpad_26
timestamp 1259953556
transform 1 0 1315 0 1 0
box -2 0 476 513
use blankpad  blankpad_25
timestamp 1259953556
transform 1 0 1789 0 1 0
box -2 0 476 513
use blankpad  blankpad_24
timestamp 1259953556
transform 1 0 2263 0 1 0
box -2 0 476 513
use blankpad  blankpad_23
timestamp 1259953556
transform 1 0 2737 0 1 0
box -2 0 476 513
use blankpad  blankpad_22
timestamp 1259953556
transform 1 0 3211 0 1 0
box -2 0 476 513
use blankpad  blankpad_21
timestamp 1259953556
transform 1 0 3685 0 1 0
box -2 0 476 513
use padframe_right  padframe_right_0
timestamp 1259953556
transform 1 0 4487 0 1 367
box 0 2 511 4264
use inorpad  inorpad_0
timestamp 1259953556
transform 0 -1 5000 1 0 367
box -2 0 476 513
use inorpad  inorpad_1
timestamp 1259953556
transform 1 0 4159 0 1 0
box -2 0 476 513
use padframe_bottom  padframe_bottom_0
timestamp 1259953556
transform 1 0 0 0 1 0
box 0 0 5000 513
<< end >>
